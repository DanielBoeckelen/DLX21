
module mux21_NBIT32_0 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n54, n59, n60, n61, n62, n63,
         n64, n65, n1, n2, n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(n7), .ZN(n2) );
  INV_X1 U2 ( .A(n7), .ZN(n1) );
  BUF_X1 U3 ( .A(n8), .Z(n5) );
  BUF_X1 U4 ( .A(n8), .Z(n6) );
  BUF_X1 U5 ( .A(n8), .Z(n3) );
  BUF_X1 U6 ( .A(n8), .Z(n4) );
  BUF_X1 U7 ( .A(n8), .Z(n7) );
  INV_X1 U8 ( .A(S), .ZN(n8) );
  INV_X1 U9 ( .A(n63), .ZN(Z[11]) );
  AOI22_X1 U10 ( .A1(A[11]), .A2(n3), .B1(B[11]), .B2(n2), .ZN(n63) );
  INV_X1 U11 ( .A(n61), .ZN(Z[13]) );
  AOI22_X1 U12 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n1), .ZN(n61) );
  INV_X1 U13 ( .A(n60), .ZN(Z[14]) );
  AOI22_X1 U14 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n1), .ZN(n60) );
  INV_X1 U15 ( .A(n54), .ZN(Z[1]) );
  AOI22_X1 U16 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n1), .ZN(n54) );
  INV_X1 U17 ( .A(n43), .ZN(Z[2]) );
  AOI22_X1 U18 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n1), .ZN(n43) );
  INV_X1 U19 ( .A(n40), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n1), .ZN(n40) );
  INV_X1 U21 ( .A(n39), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n1), .ZN(n39) );
  INV_X1 U23 ( .A(n38), .ZN(Z[5]) );
  AOI22_X1 U24 ( .A1(A[5]), .A2(n5), .B1(B[5]), .B2(n1), .ZN(n38) );
  INV_X1 U25 ( .A(n37), .ZN(Z[6]) );
  AOI22_X1 U26 ( .A1(A[6]), .A2(n6), .B1(B[6]), .B2(n1), .ZN(n37) );
  INV_X1 U27 ( .A(n35), .ZN(Z[8]) );
  AOI22_X1 U28 ( .A1(A[8]), .A2(n6), .B1(B[8]), .B2(n1), .ZN(n35) );
  INV_X1 U29 ( .A(n64), .ZN(Z[10]) );
  AOI22_X1 U30 ( .A1(A[10]), .A2(n3), .B1(B[10]), .B2(n2), .ZN(n64) );
  INV_X1 U31 ( .A(n62), .ZN(Z[12]) );
  AOI22_X1 U32 ( .A1(A[12]), .A2(n3), .B1(B[12]), .B2(n1), .ZN(n62) );
  INV_X1 U33 ( .A(n34), .ZN(Z[9]) );
  AOI22_X1 U34 ( .A1(A[9]), .A2(n6), .B1(n2), .B2(B[9]), .ZN(n34) );
  INV_X1 U35 ( .A(n65), .ZN(Z[0]) );
  AOI22_X1 U36 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n2), .ZN(n65) );
  INV_X1 U37 ( .A(n59), .ZN(Z[15]) );
  AOI22_X1 U38 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n1), .ZN(n59) );
  INV_X1 U39 ( .A(n36), .ZN(Z[7]) );
  AOI22_X1 U40 ( .A1(A[7]), .A2(n6), .B1(B[7]), .B2(n1), .ZN(n36) );
  MUX2_X1 U41 ( .A(A[16]), .B(B[16]), .S(n2), .Z(Z[16]) );
  MUX2_X1 U42 ( .A(A[17]), .B(B[17]), .S(n2), .Z(Z[17]) );
  MUX2_X1 U43 ( .A(A[18]), .B(B[18]), .S(n1), .Z(Z[18]) );
  MUX2_X1 U44 ( .A(A[19]), .B(B[19]), .S(S), .Z(Z[19]) );
  MUX2_X1 U45 ( .A(A[20]), .B(B[20]), .S(S), .Z(Z[20]) );
  MUX2_X1 U46 ( .A(A[21]), .B(B[21]), .S(S), .Z(Z[21]) );
  MUX2_X1 U47 ( .A(A[22]), .B(B[22]), .S(n2), .Z(Z[22]) );
  MUX2_X1 U48 ( .A(A[23]), .B(B[23]), .S(n2), .Z(Z[23]) );
  MUX2_X1 U49 ( .A(A[24]), .B(B[24]), .S(n2), .Z(Z[24]) );
  MUX2_X1 U50 ( .A(A[25]), .B(B[25]), .S(n2), .Z(Z[25]) );
  MUX2_X1 U51 ( .A(A[26]), .B(B[26]), .S(n2), .Z(Z[26]) );
  MUX2_X1 U52 ( .A(A[27]), .B(B[27]), .S(n2), .Z(Z[27]) );
  MUX2_X1 U53 ( .A(A[28]), .B(B[28]), .S(n2), .Z(Z[28]) );
  MUX2_X1 U54 ( .A(A[29]), .B(B[29]), .S(n2), .Z(Z[29]) );
  MUX2_X1 U55 ( .A(A[30]), .B(B[30]), .S(n2), .Z(Z[30]) );
  MUX2_X1 U56 ( .A(A[31]), .B(B[31]), .S(n2), .Z(Z[31]) );
endmodule


module mux21_NBIT32_6 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111;

  INV_X1 U1 ( .A(n15), .ZN(n5) );
  INV_X1 U2 ( .A(n15), .ZN(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n13) );
  BUF_X1 U4 ( .A(n2), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n10) );
  BUF_X1 U6 ( .A(n1), .Z(n9) );
  BUF_X1 U7 ( .A(n2), .Z(n11) );
  BUF_X1 U8 ( .A(n3), .Z(n15) );
  BUF_X1 U9 ( .A(n3), .Z(n14) );
  BUF_X1 U10 ( .A(n1), .Z(n8) );
  BUF_X1 U11 ( .A(n1), .Z(n7) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n104), .ZN(Z[31]) );
  INV_X1 U16 ( .A(n105), .ZN(Z[3]) );
  INV_X1 U17 ( .A(n106), .ZN(Z[4]) );
  INV_X1 U18 ( .A(n107), .ZN(Z[5]) );
  INV_X1 U19 ( .A(n108), .ZN(Z[6]) );
  INV_X1 U20 ( .A(n110), .ZN(Z[8]) );
  INV_X1 U21 ( .A(n81), .ZN(Z[10]) );
  INV_X1 U22 ( .A(n109), .ZN(Z[7]) );
  INV_X1 U23 ( .A(n102), .ZN(Z[2]) );
  AOI22_X1 U24 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n8), .ZN(n102) );
  INV_X1 U25 ( .A(n82), .ZN(Z[11]) );
  AOI22_X1 U26 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n14), .ZN(n82) );
  INV_X1 U27 ( .A(n83), .ZN(Z[12]) );
  AOI22_X1 U28 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n13), .ZN(n83) );
  INV_X1 U29 ( .A(n84), .ZN(Z[13]) );
  AOI22_X1 U30 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n13), .ZN(n84) );
  INV_X1 U31 ( .A(n85), .ZN(Z[14]) );
  AOI22_X1 U32 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n13), .ZN(n85) );
  INV_X1 U33 ( .A(n86), .ZN(Z[15]) );
  AOI22_X1 U34 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n13), .ZN(n86) );
  INV_X1 U35 ( .A(n87), .ZN(Z[16]) );
  AOI22_X1 U36 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n12), .ZN(n87) );
  INV_X1 U37 ( .A(n88), .ZN(Z[17]) );
  AOI22_X1 U38 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n12), .ZN(n88) );
  INV_X1 U39 ( .A(n89), .ZN(Z[18]) );
  AOI22_X1 U40 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n12), .ZN(n89) );
  INV_X1 U41 ( .A(n90), .ZN(Z[19]) );
  AOI22_X1 U42 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n12), .ZN(n90) );
  INV_X1 U43 ( .A(n92), .ZN(Z[20]) );
  AOI22_X1 U44 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n11), .ZN(n92) );
  INV_X1 U45 ( .A(n93), .ZN(Z[21]) );
  AOI22_X1 U46 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n11), .ZN(n93) );
  INV_X1 U47 ( .A(n94), .ZN(Z[22]) );
  AOI22_X1 U48 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n10), .ZN(n94) );
  INV_X1 U49 ( .A(n95), .ZN(Z[23]) );
  AOI22_X1 U50 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n10), .ZN(n95) );
  INV_X1 U51 ( .A(n96), .ZN(Z[24]) );
  AOI22_X1 U52 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n10), .ZN(n96) );
  INV_X1 U53 ( .A(n97), .ZN(Z[25]) );
  AOI22_X1 U54 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n10), .ZN(n97) );
  INV_X1 U55 ( .A(n98), .ZN(Z[26]) );
  AOI22_X1 U56 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n9), .ZN(n98) );
  INV_X1 U57 ( .A(n99), .ZN(Z[27]) );
  AOI22_X1 U58 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n9), .ZN(n99) );
  INV_X1 U59 ( .A(n100), .ZN(Z[28]) );
  AOI22_X1 U60 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n9), .ZN(n100) );
  INV_X1 U61 ( .A(n101), .ZN(Z[29]) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n9), .ZN(n101) );
  INV_X1 U63 ( .A(n103), .ZN(Z[30]) );
  AOI22_X1 U64 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n11), .ZN(n103) );
  INV_X1 U65 ( .A(n91), .ZN(Z[1]) );
  AOI22_X1 U66 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n11), .ZN(n91) );
  INV_X1 U67 ( .A(n80), .ZN(Z[0]) );
  AOI22_X1 U68 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n14), .ZN(n80) );
  INV_X1 U69 ( .A(n111), .ZN(Z[9]) );
  AOI22_X1 U70 ( .A1(A[31]), .A2(n6), .B1(B[31]), .B2(n8), .ZN(n104) );
  AOI22_X1 U71 ( .A1(A[3]), .A2(n6), .B1(B[3]), .B2(n8), .ZN(n105) );
  AOI22_X1 U72 ( .A1(A[6]), .A2(n6), .B1(B[6]), .B2(n7), .ZN(n108) );
  AOI22_X1 U73 ( .A1(A[4]), .A2(n6), .B1(B[4]), .B2(n8), .ZN(n106) );
  AOI22_X1 U74 ( .A1(A[7]), .A2(n6), .B1(B[7]), .B2(n7), .ZN(n109) );
  AOI22_X1 U75 ( .A1(A[5]), .A2(n6), .B1(B[5]), .B2(n7), .ZN(n107) );
  AOI22_X1 U76 ( .A1(A[9]), .A2(n6), .B1(n14), .B2(B[9]), .ZN(n111) );
  AOI22_X1 U77 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n14), .ZN(n81) );
  AOI22_X1 U78 ( .A1(A[8]), .A2(n6), .B1(B[8]), .B2(n7), .ZN(n110) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module mux21_NBIT32_5 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n3), .Z(n14) );
  BUF_X1 U8 ( .A(n3), .Z(n13) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n2), .Z(n10) );
  BUF_X1 U11 ( .A(n1), .Z(n8) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n1) );
  BUF_X1 U14 ( .A(S), .Z(n2) );
  INV_X1 U15 ( .A(n98), .ZN(Z[27]) );
  INV_X1 U16 ( .A(n97), .ZN(Z[26]) );
  INV_X1 U17 ( .A(n100), .ZN(Z[29]) );
  INV_X1 U18 ( .A(n102), .ZN(Z[30]) );
  INV_X1 U19 ( .A(n103), .ZN(Z[31]) );
  INV_X1 U20 ( .A(n99), .ZN(Z[28]) );
  INV_X1 U21 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U22 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U23 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U24 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U25 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U26 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U27 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U28 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U29 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U30 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U31 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U32 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U33 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U34 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U35 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U36 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U37 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U38 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U39 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U40 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U41 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U42 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U43 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U44 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U45 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U46 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U47 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U48 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U49 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U50 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U51 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U52 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U53 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U54 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U55 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U56 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U57 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U58 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U59 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U60 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U61 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U62 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U63 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U64 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U65 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U66 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U67 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U68 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U69 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U70 ( .A1(A[9]), .A2(n4), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U71 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U72 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  AOI22_X1 U73 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  AOI22_X1 U74 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  AOI22_X1 U75 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  AOI22_X1 U76 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  AOI22_X1 U77 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n5), .B1(B[31]), .B2(n7), .ZN(n103) );
endmodule


module regn_N32_0 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n17, n18, n19;

  DFFR_X1 DOUT_reg_31_ ( .D(n96), .CK(CLK), .RN(n19), .Q(DOUT[31]) );
  DFFR_X1 DOUT_reg_30_ ( .D(n95), .CK(CLK), .RN(n19), .Q(DOUT[30]) );
  DFFR_X1 DOUT_reg_29_ ( .D(n94), .CK(CLK), .RN(n19), .Q(DOUT[29]) );
  DFFR_X1 DOUT_reg_28_ ( .D(n93), .CK(CLK), .RN(n19), .Q(DOUT[28]) );
  DFFR_X1 DOUT_reg_27_ ( .D(n92), .CK(CLK), .RN(n19), .Q(DOUT[27]) );
  DFFR_X1 DOUT_reg_26_ ( .D(n91), .CK(CLK), .RN(n19), .Q(DOUT[26]) );
  DFFR_X1 DOUT_reg_25_ ( .D(n90), .CK(CLK), .RN(n19), .Q(DOUT[25]) );
  DFFR_X1 DOUT_reg_24_ ( .D(n89), .CK(CLK), .RN(n19), .Q(DOUT[24]) );
  DFFR_X1 DOUT_reg_23_ ( .D(n88), .CK(CLK), .RN(n18), .Q(DOUT[23]) );
  DFFR_X1 DOUT_reg_22_ ( .D(n87), .CK(CLK), .RN(n18), .Q(DOUT[22]) );
  DFFR_X1 DOUT_reg_21_ ( .D(n86), .CK(CLK), .RN(n18), .Q(DOUT[21]) );
  DFFR_X1 DOUT_reg_20_ ( .D(n85), .CK(CLK), .RN(n18), .Q(DOUT[20]) );
  DFFR_X1 DOUT_reg_19_ ( .D(n84), .CK(CLK), .RN(n18), .Q(DOUT[19]) );
  DFFR_X1 DOUT_reg_18_ ( .D(n83), .CK(CLK), .RN(n18), .Q(DOUT[18]) );
  DFFR_X1 DOUT_reg_17_ ( .D(n82), .CK(CLK), .RN(n18), .Q(DOUT[17]) );
  DFFR_X1 DOUT_reg_16_ ( .D(n81), .CK(CLK), .RN(n18), .Q(DOUT[16]) );
  DFFR_X1 DOUT_reg_15_ ( .D(n80), .CK(CLK), .RN(n18), .Q(DOUT[15]), .QN(n48)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n79), .CK(CLK), .RN(n18), .Q(DOUT[14]), .QN(n47)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n78), .CK(CLK), .RN(n18), .Q(DOUT[13]), .QN(n46)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n77), .CK(CLK), .RN(n18), .Q(DOUT[12]), .QN(n45)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n76), .CK(CLK), .RN(n17), .Q(DOUT[11]), .QN(n44)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n75), .CK(CLK), .RN(n17), .Q(DOUT[10]), .QN(n43)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n74), .CK(CLK), .RN(n17), .Q(DOUT[9]), .QN(n42) );
  DFFR_X1 DOUT_reg_8_ ( .D(n73), .CK(CLK), .RN(n17), .Q(DOUT[8]), .QN(n41) );
  DFFR_X1 DOUT_reg_7_ ( .D(n72), .CK(CLK), .RN(n17), .Q(DOUT[7]), .QN(n40) );
  DFFR_X1 DOUT_reg_6_ ( .D(n71), .CK(CLK), .RN(n17), .Q(DOUT[6]), .QN(n39) );
  DFFR_X1 DOUT_reg_5_ ( .D(n70), .CK(CLK), .RN(n17), .Q(DOUT[5]), .QN(n38) );
  DFFR_X1 DOUT_reg_4_ ( .D(n69), .CK(CLK), .RN(n17), .Q(DOUT[4]), .QN(n37) );
  DFFR_X1 DOUT_reg_3_ ( .D(n68), .CK(CLK), .RN(n17), .Q(DOUT[3]), .QN(n36) );
  DFFR_X1 DOUT_reg_2_ ( .D(n67), .CK(CLK), .RN(n17), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 DOUT_reg_1_ ( .D(n66), .CK(CLK), .RN(n17), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 DOUT_reg_0_ ( .D(n65), .CK(CLK), .RN(n17), .Q(DOUT[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RST), .Z(n17) );
  BUF_X1 U3 ( .A(RST), .Z(n18) );
  BUF_X1 U4 ( .A(RST), .Z(n19) );
  OAI21_X1 U5 ( .B1(n44), .B2(EN), .A(n12), .ZN(n76) );
  NAND2_X1 U6 ( .A1(DIN[11]), .A2(EN), .ZN(n12) );
  OAI21_X1 U7 ( .B1(n46), .B2(EN), .A(n14), .ZN(n78) );
  NAND2_X1 U8 ( .A1(DIN[13]), .A2(EN), .ZN(n14) );
  OAI21_X1 U9 ( .B1(n47), .B2(EN), .A(n15), .ZN(n79) );
  NAND2_X1 U10 ( .A1(DIN[14]), .A2(EN), .ZN(n15) );
  OAI21_X1 U11 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U12 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U13 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U14 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U15 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U16 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U17 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X1 U18 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U19 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X1 U20 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U21 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U22 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X1 U23 ( .B1(n41), .B2(EN), .A(n9), .ZN(n73) );
  NAND2_X1 U24 ( .A1(DIN[8]), .A2(EN), .ZN(n9) );
  OAI21_X1 U25 ( .B1(n43), .B2(EN), .A(n11), .ZN(n75) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n11) );
  OAI21_X1 U27 ( .B1(n45), .B2(EN), .A(n13), .ZN(n77) );
  NAND2_X1 U28 ( .A1(DIN[12]), .A2(EN), .ZN(n13) );
  OAI21_X1 U29 ( .B1(n42), .B2(EN), .A(n10), .ZN(n74) );
  NAND2_X1 U30 ( .A1(DIN[9]), .A2(EN), .ZN(n10) );
  OAI21_X1 U31 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U32 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U33 ( .B1(n48), .B2(EN), .A(n16), .ZN(n80) );
  NAND2_X1 U34 ( .A1(DIN[15]), .A2(EN), .ZN(n16) );
  NAND2_X1 U35 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X1 U36 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  MUX2_X1 U37 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n81) );
  MUX2_X1 U38 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n82) );
  MUX2_X1 U39 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n83) );
  MUX2_X1 U40 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n84) );
  MUX2_X1 U41 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U42 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U43 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U44 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n88) );
  MUX2_X1 U45 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U46 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n90) );
  MUX2_X1 U47 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U48 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n92) );
  MUX2_X1 U49 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n93) );
  MUX2_X1 U50 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n94) );
  MUX2_X1 U51 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
  MUX2_X1 U52 ( .A(DOUT[31]), .B(DIN[31]), .S(EN), .Z(n96) );
endmodule


module regn_N32_9 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U6 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U7 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U8 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U9 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U10 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U11 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U12 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U13 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U14 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U15 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U16 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U17 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U18 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U22 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U23 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U24 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U25 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U26 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U27 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U28 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U29 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U30 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U31 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U32 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U33 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U34 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U35 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U36 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U37 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U38 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U39 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U40 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U41 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U42 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U43 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U44 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U45 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U46 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U47 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U48 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U49 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U50 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U51 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U52 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U53 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U54 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U55 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U56 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U57 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U58 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U59 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U60 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U61 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U62 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U63 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U64 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U65 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U66 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U67 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U68 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
endmodule


module regn_N32_8 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197;

  DFFR_X1 DOUT_reg_25_ ( .D(n108), .CK(CLK), .RN(n101), .Q(DOUT[25]), .QN(n140) );
  DFFR_X1 DOUT_reg_24_ ( .D(n109), .CK(CLK), .RN(n101), .Q(DOUT[24]), .QN(n141) );
  DFFR_X1 DOUT_reg_23_ ( .D(n110), .CK(CLK), .RN(n100), .Q(DOUT[23]), .QN(n142) );
  DFFR_X1 DOUT_reg_22_ ( .D(n111), .CK(CLK), .RN(n100), .Q(DOUT[22]), .QN(n143) );
  DFFR_X1 DOUT_reg_21_ ( .D(n112), .CK(CLK), .RN(n100), .Q(DOUT[21]), .QN(n144) );
  DFFR_X1 DOUT_reg_20_ ( .D(n113), .CK(CLK), .RN(n100), .Q(DOUT[20]), .QN(n145) );
  DFFR_X1 DOUT_reg_19_ ( .D(n114), .CK(CLK), .RN(n100), .Q(DOUT[19]), .QN(n146) );
  DFFR_X1 DOUT_reg_18_ ( .D(n115), .CK(CLK), .RN(n100), .Q(DOUT[18]), .QN(n147) );
  DFFR_X1 DOUT_reg_17_ ( .D(n116), .CK(CLK), .RN(n100), .Q(DOUT[17]), .QN(n148) );
  DFFR_X1 DOUT_reg_16_ ( .D(n117), .CK(CLK), .RN(n100), .Q(DOUT[16]), .QN(n149) );
  DFFR_X1 DOUT_reg_15_ ( .D(n118), .CK(CLK), .RN(n100), .Q(DOUT[15]), .QN(n150) );
  DFFR_X1 DOUT_reg_14_ ( .D(n119), .CK(CLK), .RN(n100), .Q(DOUT[14]), .QN(n151) );
  DFFR_X1 DOUT_reg_13_ ( .D(n120), .CK(CLK), .RN(n100), .Q(DOUT[13]), .QN(n152) );
  DFFR_X1 DOUT_reg_12_ ( .D(n121), .CK(CLK), .RN(n100), .Q(DOUT[12]), .QN(n153) );
  DFFR_X1 DOUT_reg_11_ ( .D(n122), .CK(CLK), .RN(n99), .Q(DOUT[11]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n123), .CK(CLK), .RN(n99), .Q(DOUT[10]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n124), .CK(CLK), .RN(n99), .Q(DOUT[9]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n125), .CK(CLK), .RN(n99), .Q(DOUT[8]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n126), .CK(CLK), .RN(n99), .Q(DOUT[7]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n127), .CK(CLK), .RN(n99), .Q(DOUT[6]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n128), .CK(CLK), .RN(n99), .Q(DOUT[5]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n129), .CK(CLK), .RN(n99), .Q(DOUT[4]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n130), .CK(CLK), .RN(n99), .Q(DOUT[3]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n131), .CK(CLK), .RN(n99), .Q(DOUT[2]), .QN(n163)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n132), .CK(CLK), .RN(n99), .Q(DOUT[1]), .QN(n164)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n133), .CK(CLK), .RN(n99), .Q(DOUT[0]), .QN(n165)
         );
  DFFR_X1 DOUT_reg_31_ ( .D(n102), .CK(CLK), .RN(n101), .Q(DOUT[31]), .QN(n134) );
  DFFR_X1 DOUT_reg_28_ ( .D(n105), .CK(CLK), .RN(n101), .QN(n137) );
  DFFR_X1 DOUT_reg_30_ ( .D(n103), .CK(CLK), .RN(n101), .Q(DOUT[30]), .QN(n135) );
  DFFR_X1 DOUT_reg_29_ ( .D(n104), .CK(CLK), .RN(n101), .Q(DOUT[29]), .QN(n136) );
  DFFR_X1 DOUT_reg_26_ ( .D(n107), .CK(CLK), .RN(n101), .Q(DOUT[26]), .QN(n139) );
  DFFR_X1 DOUT_reg_27_ ( .D(n106), .CK(CLK), .RN(n101), .Q(DOUT[27]), .QN(n138) );
  INV_X2 U2 ( .A(n137), .ZN(DOUT[28]) );
  BUF_X1 U3 ( .A(RST), .Z(n99) );
  BUF_X1 U4 ( .A(RST), .Z(n100) );
  BUF_X1 U5 ( .A(RST), .Z(n101) );
  NAND2_X1 U6 ( .A1(DIN[27]), .A2(EN), .ZN(n170) );
  NAND2_X1 U7 ( .A1(DIN[26]), .A2(EN), .ZN(n171) );
  NAND2_X1 U8 ( .A1(DIN[29]), .A2(EN), .ZN(n168) );
  NAND2_X1 U9 ( .A1(DIN[30]), .A2(EN), .ZN(n167) );
  NAND2_X1 U10 ( .A1(DIN[31]), .A2(EN), .ZN(n166) );
  NAND2_X1 U11 ( .A1(DIN[28]), .A2(EN), .ZN(n169) );
  OAI21_X1 U12 ( .B1(n164), .B2(EN), .A(n196), .ZN(n132) );
  NAND2_X1 U13 ( .A1(DIN[1]), .A2(EN), .ZN(n196) );
  OAI21_X1 U14 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U15 ( .A1(DIN[2]), .A2(EN), .ZN(n195) );
  OAI21_X1 U16 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U17 ( .A1(DIN[3]), .A2(EN), .ZN(n194) );
  OAI21_X1 U18 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U19 ( .A1(DIN[4]), .A2(EN), .ZN(n193) );
  OAI21_X1 U20 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U21 ( .A1(DIN[5]), .A2(EN), .ZN(n192) );
  OAI21_X1 U22 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U23 ( .A1(DIN[6]), .A2(EN), .ZN(n191) );
  OAI21_X1 U24 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U25 ( .A1(DIN[7]), .A2(EN), .ZN(n190) );
  OAI21_X1 U26 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U27 ( .A1(DIN[8]), .A2(EN), .ZN(n189) );
  OAI21_X1 U28 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U29 ( .A1(DIN[10]), .A2(EN), .ZN(n187) );
  OAI21_X1 U30 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U31 ( .A1(DIN[11]), .A2(EN), .ZN(n186) );
  OAI21_X1 U32 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U33 ( .A1(DIN[12]), .A2(EN), .ZN(n185) );
  OAI21_X1 U34 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U35 ( .A1(DIN[13]), .A2(EN), .ZN(n184) );
  OAI21_X1 U36 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U37 ( .A1(DIN[14]), .A2(EN), .ZN(n183) );
  OAI21_X1 U38 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U39 ( .A1(DIN[15]), .A2(EN), .ZN(n182) );
  OAI21_X1 U40 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U41 ( .A1(DIN[16]), .A2(EN), .ZN(n181) );
  OAI21_X1 U42 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U43 ( .A1(DIN[17]), .A2(EN), .ZN(n180) );
  OAI21_X1 U44 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U45 ( .A1(DIN[18]), .A2(EN), .ZN(n179) );
  OAI21_X1 U46 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U47 ( .A1(DIN[19]), .A2(EN), .ZN(n178) );
  OAI21_X1 U48 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U49 ( .A1(DIN[20]), .A2(EN), .ZN(n177) );
  OAI21_X1 U50 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U51 ( .A1(DIN[21]), .A2(EN), .ZN(n176) );
  OAI21_X1 U52 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U53 ( .A1(DIN[22]), .A2(EN), .ZN(n175) );
  OAI21_X1 U54 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U55 ( .A1(DIN[23]), .A2(EN), .ZN(n174) );
  OAI21_X1 U56 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U57 ( .A1(DIN[24]), .A2(EN), .ZN(n173) );
  OAI21_X1 U58 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U59 ( .A1(DIN[25]), .A2(EN), .ZN(n172) );
  OAI21_X1 U60 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U61 ( .A1(DIN[9]), .A2(EN), .ZN(n188) );
  OAI21_X1 U62 ( .B1(n165), .B2(EN), .A(n197), .ZN(n133) );
  NAND2_X1 U63 ( .A1(EN), .A2(DIN[0]), .ZN(n197) );
  OAI21_X1 U64 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  OAI21_X1 U65 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  OAI21_X1 U66 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  OAI21_X1 U67 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  OAI21_X1 U68 ( .B1(EN), .B2(n137), .A(n169), .ZN(n105) );
  OAI21_X1 U69 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
endmodule


module Fetch_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XOR2_X1 U2 ( .A(n1), .B(n18), .Z(SUM[31]) );
  NAND2_X1 U3 ( .A1(n19), .A2(A[30]), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n69), .A2(n52), .ZN(n13) );
  AND2_X1 U5 ( .A1(n13), .A2(n11), .ZN(n58) );
  NOR2_X1 U6 ( .A1(n70), .A2(n12), .ZN(n62) );
  INV_X1 U7 ( .A(n32), .ZN(n36) );
  INV_X1 U8 ( .A(n25), .ZN(n29) );
  INV_X1 U9 ( .A(n40), .ZN(n44) );
  OR2_X1 U10 ( .A1(n32), .A2(n33), .ZN(n2) );
  NOR2_X1 U11 ( .A1(n4), .A2(n5), .ZN(n3) );
  NAND3_X1 U12 ( .A1(n50), .A2(n51), .A3(n11), .ZN(n4) );
  OR2_X1 U13 ( .A1(n48), .A2(n49), .ZN(n5) );
  AND2_X1 U14 ( .A1(n57), .A2(A[13]), .ZN(n54) );
  AND2_X1 U15 ( .A1(n15), .A2(A[5]), .ZN(n14) );
  NOR2_X1 U16 ( .A1(n32), .A2(n33), .ZN(n30) );
  NOR2_X1 U17 ( .A1(n9), .A2(n21), .ZN(n19) );
  AND2_X1 U18 ( .A1(A[12]), .A2(n58), .ZN(n57) );
  NOR2_X1 U19 ( .A1(n68), .A2(n69), .ZN(n15) );
  NOR2_X1 U20 ( .A1(n40), .A2(n41), .ZN(n37) );
  AND4_X1 U21 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n11) );
  NOR2_X1 U22 ( .A1(n25), .A2(n26), .ZN(n23) );
  NOR2_X1 U23 ( .A1(SUM[2]), .A2(n16), .ZN(n51) );
  AND2_X1 U24 ( .A1(n54), .A2(A[14]), .ZN(n53) );
  AND2_X1 U25 ( .A1(n62), .A2(A[10]), .ZN(n61) );
  AND2_X1 U26 ( .A1(n8), .A2(A[18]), .ZN(n42) );
  NAND2_X1 U27 ( .A1(n13), .A2(A[8]), .ZN(n12) );
  AND2_X1 U28 ( .A1(A[21]), .A2(n36), .ZN(n6) );
  AND2_X1 U29 ( .A1(A[25]), .A2(n29), .ZN(n7) );
  AND2_X1 U30 ( .A1(A[17]), .A2(n44), .ZN(n8) );
  NAND2_X1 U31 ( .A1(A[22]), .A2(n6), .ZN(n34) );
  NAND2_X1 U32 ( .A1(A[26]), .A2(n7), .ZN(n27) );
  NAND2_X1 U33 ( .A1(A[12]), .A2(A[13]), .ZN(n49) );
  NAND2_X1 U34 ( .A1(A[14]), .A2(A[15]), .ZN(n48) );
  NAND2_X1 U35 ( .A1(n23), .A2(A[28]), .ZN(n9) );
  AND2_X1 U36 ( .A1(A[6]), .A2(n14), .ZN(n10) );
  INV_X1 U37 ( .A(A[14]), .ZN(n56) );
  INV_X1 U38 ( .A(A[3]), .ZN(n16) );
  INV_X1 U39 ( .A(A[29]), .ZN(n21) );
  XNOR2_X1 U40 ( .A(n65), .B(n10), .ZN(SUM[7]) );
  XNOR2_X1 U41 ( .A(n68), .B(n51), .ZN(SUM[4]) );
  INV_X1 U42 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U43 ( .A(A[13]), .ZN(n59) );
  INV_X1 U44 ( .A(A[12]), .ZN(n60) );
  INV_X1 U45 ( .A(A[17]), .ZN(n46) );
  INV_X1 U46 ( .A(A[25]), .ZN(n31) );
  INV_X1 U47 ( .A(A[26]), .ZN(n28) );
  INV_X1 U48 ( .A(A[18]), .ZN(n45) );
  INV_X1 U49 ( .A(A[15]), .ZN(n55) );
  XNOR2_X1 U50 ( .A(n66), .B(n14), .ZN(SUM[6]) );
  XNOR2_X1 U51 ( .A(n56), .B(n54), .ZN(SUM[14]) );
  XNOR2_X1 U52 ( .A(n16), .B(A[2]), .ZN(SUM[3]) );
  XNOR2_X1 U53 ( .A(n60), .B(n58), .ZN(SUM[12]) );
  XNOR2_X1 U54 ( .A(n6), .B(n35), .ZN(SUM[22]) );
  XNOR2_X1 U55 ( .A(n34), .B(A[23]), .ZN(SUM[23]) );
  XNOR2_X1 U56 ( .A(n2), .B(A[24]), .ZN(SUM[24]) );
  XNOR2_X1 U57 ( .A(n31), .B(n29), .ZN(SUM[25]) );
  XNOR2_X1 U58 ( .A(n7), .B(n28), .ZN(SUM[26]) );
  XNOR2_X1 U59 ( .A(n24), .B(A[28]), .ZN(SUM[28]) );
  XNOR2_X1 U60 ( .A(n21), .B(n22), .ZN(SUM[29]) );
  XNOR2_X1 U61 ( .A(n27), .B(A[27]), .ZN(SUM[27]) );
  XNOR2_X1 U62 ( .A(n38), .B(n36), .ZN(SUM[21]) );
  XNOR2_X1 U63 ( .A(n45), .B(n8), .ZN(SUM[18]) );
  XNOR2_X1 U64 ( .A(n46), .B(n44), .ZN(SUM[17]) );
  INV_X1 U65 ( .A(A[19]), .ZN(n43) );
  INV_X1 U66 ( .A(A[11]), .ZN(n63) );
  INV_X1 U67 ( .A(A[21]), .ZN(n38) );
  INV_X1 U68 ( .A(A[22]), .ZN(n35) );
  INV_X1 U69 ( .A(A[31]), .ZN(n18) );
  INV_X1 U70 ( .A(A[6]), .ZN(n66) );
  INV_X1 U71 ( .A(A[4]), .ZN(n68) );
  INV_X1 U72 ( .A(n9), .ZN(n22) );
  INV_X1 U73 ( .A(A[7]), .ZN(n65) );
  INV_X1 U74 ( .A(A[5]), .ZN(n67) );
  INV_X1 U75 ( .A(A[9]), .ZN(n70) );
  INV_X1 U76 ( .A(A[10]), .ZN(n71) );
  NAND4_X1 U77 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n52) );
  NAND2_X1 U78 ( .A1(n37), .A2(A[20]), .ZN(n32) );
  NAND2_X1 U79 ( .A1(n30), .A2(A[24]), .ZN(n25) );
  NAND2_X1 U80 ( .A1(n3), .A2(A[16]), .ZN(n40) );
  XNOR2_X1 U81 ( .A(n20), .B(A[30]), .ZN(SUM[30]) );
  INV_X1 U82 ( .A(A[8]), .ZN(n64) );
  XNOR2_X1 U83 ( .A(n12), .B(A[9]), .ZN(SUM[9]) );
  XNOR2_X1 U84 ( .A(n64), .B(n13), .ZN(SUM[8]) );
  XNOR2_X1 U85 ( .A(n67), .B(n15), .ZN(SUM[5]) );
  INV_X1 U86 ( .A(n19), .ZN(n20) );
  INV_X1 U87 ( .A(n23), .ZN(n24) );
  NAND3_X1 U88 ( .A1(A[26]), .A2(A[27]), .A3(A[25]), .ZN(n26) );
  NAND3_X1 U89 ( .A1(A[22]), .A2(A[23]), .A3(A[21]), .ZN(n33) );
  XNOR2_X1 U90 ( .A(n39), .B(A[20]), .ZN(SUM[20]) );
  INV_X1 U91 ( .A(n37), .ZN(n39) );
  NAND3_X1 U92 ( .A1(A[18]), .A2(A[19]), .A3(A[17]), .ZN(n41) );
  XNOR2_X1 U93 ( .A(n43), .B(n42), .ZN(SUM[19]) );
  XNOR2_X1 U94 ( .A(n47), .B(A[16]), .ZN(SUM[16]) );
  INV_X1 U95 ( .A(n3), .ZN(n47) );
  INV_X1 U96 ( .A(n52), .ZN(n50) );
  XNOR2_X1 U97 ( .A(n55), .B(n53), .ZN(SUM[15]) );
  XNOR2_X1 U98 ( .A(n59), .B(n57), .ZN(SUM[13]) );
  XNOR2_X1 U99 ( .A(n63), .B(n61), .ZN(SUM[11]) );
  XNOR2_X1 U100 ( .A(n71), .B(n62), .ZN(SUM[10]) );
  INV_X1 U101 ( .A(n51), .ZN(n69) );
endmodule


module Fetch ( CLK, RST, ZERO_FLAG, PC_EXT, INS_IN, Bubble_in, HDU_INS_IN, 
        HDU_PC_IN, HDU_NPC_IN, PC_OUT, ADDR_OUT, NPC_OUT, INS_OUT );
  input [31:0] PC_EXT;
  input [31:0] INS_IN;
  input [31:0] HDU_INS_IN;
  input [31:0] HDU_PC_IN;
  input [31:0] HDU_NPC_IN;
  output [31:0] PC_OUT;
  output [31:0] ADDR_OUT;
  output [31:0] NPC_OUT;
  output [31:0] INS_OUT;
  input CLK, RST, ZERO_FLAG, Bubble_in;
  wire   n6, sig_RST, n5;
  wire   [31:0] sig_NPC;
  wire   [31:0] PC_MUX_OUT;
  wire   [31:0] sig_INS;

  mux21_NBIT32_0 NPC_or_NPC_HDU ( .A(PC_EXT), .B(HDU_NPC_IN), .S(Bubble_in), 
        .Z(sig_NPC) );
  mux21_NBIT32_6 PC_or_PC_HDU ( .A(ADDR_OUT), .B(HDU_PC_IN), .S(Bubble_in), 
        .Z(PC_MUX_OUT) );
  mux21_NBIT32_5 INS_or_HDU_INS ( .A(INS_IN), .B(HDU_INS_IN), .S(Bubble_in), 
        .Z(sig_INS) );
  regn_N32_0 PC ( .DIN(sig_NPC), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT({
        ADDR_OUT[31:8], n6, ADDR_OUT[6:0]}) );
  regn_N32_9 PC_reg ( .DIN(PC_MUX_OUT), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(PC_OUT) );
  regn_N32_8 IR ( .DIN(sig_INS), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        INS_OUT) );
  Fetch_DW01_add_1 add_54 ( .A({ADDR_OUT[31:8], n6, ADDR_OUT[6:0]}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC_OUT)
         );
  NOR2_X1 U6 ( .A1(ZERO_FLAG), .A2(n5), .ZN(sig_RST) );
  CLKBUF_X1 U7 ( .A(n6), .Z(ADDR_OUT[7]) );
  INV_X1 U8 ( .A(RST), .ZN(n5) );
endmodule


module instruction_type ( INST_IN, Rtype, Itype, Jtype );
  input [31:0] INST_IN;
  output Rtype, Itype, Jtype;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n1, n2, n3, n4, n5, n6, n22, n23, n24, n25, n26, n27, n28;

  OAI33_X1 U24 ( .A1(n15), .A2(n25), .A3(n11), .B1(n16), .B2(n1), .B3(
        INST_IN[28]), .ZN(n14) );
  INV_X1 U1 ( .A(n17), .ZN(n23) );
  NOR2_X1 U2 ( .A1(n7), .A2(n28), .ZN(Rtype) );
  NOR2_X1 U3 ( .A1(n27), .A2(n7), .ZN(Jtype) );
  INV_X1 U4 ( .A(n25), .ZN(n1) );
  NOR2_X1 U5 ( .A1(INST_IN[27]), .A2(INST_IN[26]), .ZN(n2) );
  NOR2_X1 U6 ( .A1(INST_IN[27]), .A2(INST_IN[26]), .ZN(n8) );
  OR2_X1 U7 ( .A1(n9), .A2(n27), .ZN(n3) );
  OR2_X1 U8 ( .A1(n10), .A2(n11), .ZN(n4) );
  NAND3_X1 U9 ( .A1(n12), .A2(n4), .A3(n3), .ZN(Itype) );
  OR2_X1 U10 ( .A1(INST_IN[29]), .A2(INST_IN[30]), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n5), .A2(n20), .ZN(n18) );
  CLKBUF_X1 U12 ( .A(INST_IN[31]), .Z(n6) );
  INV_X1 U13 ( .A(n2), .ZN(n28) );
  INV_X1 U14 ( .A(INST_IN[29]), .ZN(n26) );
  NAND2_X1 U15 ( .A1(INST_IN[26]), .A2(n27), .ZN(n11) );
  INV_X1 U16 ( .A(INST_IN[30]), .ZN(n25) );
  AOI21_X1 U17 ( .B1(INST_IN[26]), .B2(INST_IN[27]), .A(n8), .ZN(n16) );
  INV_X1 U18 ( .A(INST_IN[27]), .ZN(n27) );
  AND2_X1 U19 ( .A1(INST_IN[28]), .A2(INST_IN[30]), .ZN(n22) );
  NOR2_X1 U20 ( .A1(n22), .A2(n20), .ZN(n19) );
  NAND2_X1 U21 ( .A1(INST_IN[29]), .A2(INST_IN[28]), .ZN(n15) );
  NAND4_X1 U22 ( .A1(INST_IN[30]), .A2(INST_IN[28]), .A3(n26), .A4(n24), .ZN(
        n17) );
  NAND2_X1 U23 ( .A1(n24), .A2(INST_IN[29]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(n10), .A2(n17), .ZN(n13) );
  NOR3_X1 U26 ( .A1(n21), .A2(n23), .A3(n19), .ZN(n9) );
  AOI211_X1 U27 ( .C1(n6), .C2(n26), .A(n25), .B(INST_IN[28]), .ZN(n21) );
  OR4_X1 U28 ( .A1(INST_IN[28]), .A2(INST_IN[29]), .A3(n1), .A4(INST_IN[31]), 
        .ZN(n7) );
  AOI21_X1 U29 ( .B1(INST_IN[28]), .B2(n18), .A(n19), .ZN(n10) );
  INV_X1 U30 ( .A(INST_IN[31]), .ZN(n24) );
  AOI22_X1 U31 ( .A1(n13), .A2(n2), .B1(n6), .B2(n14), .ZN(n12) );
endmodule


module instruction_decomposition ( INST_IN, Rtype, Itype, Jtype, ADD_RS1, 
        ADD_RS2, ADD_WR, IMM, RD1, RD2 );
  input [31:0] INST_IN;
  output [4:0] ADD_RS1;
  output [4:0] ADD_RS2;
  output [4:0] ADD_WR;
  output [31:0] IMM;
  input Rtype, Itype, Jtype;
  output RD1, RD2;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n1,
         n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n38, n39, n40, n41, n42;
  assign IMM[25] = IMM[31];
  assign IMM[26] = IMM[31];
  assign IMM[27] = IMM[31];
  assign IMM[28] = IMM[31];
  assign IMM[29] = IMM[31];
  assign IMM[30] = IMM[31];

  NOR2_X2 U42 ( .A1(n5), .A2(n20), .ZN(ADD_RS2[4]) );
  NOR2_X2 U44 ( .A1(n6), .A2(n22), .ZN(ADD_RS2[2]) );
  NOR2_X2 U46 ( .A1(n3), .A2(n24), .ZN(ADD_RS2[0]) );
  NOR2_X2 U54 ( .A1(n4), .A2(n19), .ZN(ADD_RS1[0]) );
  NAND3_X1 U80 ( .A1(n11), .A2(INST_IN[26]), .A3(INST_IN[30]), .ZN(n34) );
  XOR2_X1 U81 ( .A(INST_IN[26]), .B(n15), .Z(n36) );
  AND2_X1 U3 ( .A1(n2), .A2(INST_IN[22]), .ZN(ADD_RS1[1]) );
  AND2_X1 U4 ( .A1(n2), .A2(INST_IN[24]), .ZN(ADD_RS1[3]) );
  AND2_X1 U5 ( .A1(n2), .A2(INST_IN[25]), .ZN(ADD_RS1[4]) );
  AND2_X2 U6 ( .A1(n13), .A2(n35), .ZN(n3) );
  CLKBUF_X1 U7 ( .A(Itype), .Z(n1) );
  AND2_X1 U8 ( .A1(RD1), .A2(INST_IN[23]), .ZN(ADD_RS1[2]) );
  OR2_X1 U9 ( .A1(Rtype), .A2(Itype), .ZN(n2) );
  OR2_X1 U10 ( .A1(Rtype), .A2(Itype), .ZN(RD1) );
  AND2_X1 U11 ( .A1(n13), .A2(n35), .ZN(n5) );
  INV_X1 U12 ( .A(n30), .ZN(n12) );
  INV_X1 U13 ( .A(n31), .ZN(n11) );
  INV_X1 U14 ( .A(Rtype), .ZN(n13) );
  OAI221_X1 U15 ( .B1(n31), .B2(n24), .C1(n42), .C2(n13), .A(n7), .ZN(
        ADD_WR[0]) );
  OAI221_X1 U16 ( .B1(n31), .B2(n23), .C1(n41), .C2(n13), .A(n7), .ZN(
        ADD_WR[1]) );
  OAI221_X1 U17 ( .B1(n31), .B2(n22), .C1(n40), .C2(n13), .A(n7), .ZN(
        ADD_WR[2]) );
  OAI221_X1 U18 ( .B1(n31), .B2(n21), .C1(n39), .C2(n13), .A(n7), .ZN(
        ADD_WR[3]) );
  OAI221_X1 U19 ( .B1(n31), .B2(n20), .C1(n38), .C2(n13), .A(n7), .ZN(
        ADD_WR[4]) );
  NAND2_X1 U20 ( .A1(n11), .A2(INST_IN[15]), .ZN(n29) );
  INV_X1 U21 ( .A(n25), .ZN(IMM[31]) );
  OAI21_X1 U22 ( .B1(n26), .B2(n27), .A(n13), .ZN(n25) );
  INV_X1 U23 ( .A(n32), .ZN(n7) );
  OAI21_X1 U24 ( .B1(n33), .B2(n34), .A(n28), .ZN(n32) );
  INV_X1 U25 ( .A(INST_IN[16]), .ZN(n24) );
  INV_X1 U26 ( .A(INST_IN[20]), .ZN(n20) );
  INV_X1 U27 ( .A(INST_IN[18]), .ZN(n22) );
  INV_X1 U28 ( .A(INST_IN[15]), .ZN(n38) );
  INV_X1 U29 ( .A(INST_IN[19]), .ZN(n21) );
  INV_X1 U30 ( .A(INST_IN[17]), .ZN(n23) );
  INV_X1 U31 ( .A(INST_IN[21]), .ZN(n19) );
  INV_X1 U32 ( .A(INST_IN[11]), .ZN(n42) );
  INV_X1 U33 ( .A(INST_IN[12]), .ZN(n41) );
  INV_X1 U34 ( .A(INST_IN[13]), .ZN(n40) );
  INV_X1 U35 ( .A(INST_IN[14]), .ZN(n39) );
  OAI21_X1 U36 ( .B1(n28), .B2(n24), .A(n29), .ZN(IMM[16]) );
  OAI21_X1 U37 ( .B1(n28), .B2(n23), .A(n29), .ZN(IMM[17]) );
  OAI21_X1 U38 ( .B1(n28), .B2(n22), .A(n29), .ZN(IMM[18]) );
  OAI21_X1 U39 ( .B1(n28), .B2(n21), .A(n29), .ZN(IMM[19]) );
  OAI21_X1 U40 ( .B1(n28), .B2(n20), .A(n29), .ZN(IMM[20]) );
  OAI21_X1 U41 ( .B1(n28), .B2(n19), .A(n29), .ZN(IMM[21]) );
  OAI21_X1 U43 ( .B1(n28), .B2(n18), .A(n29), .ZN(IMM[22]) );
  OAI21_X1 U45 ( .B1(n28), .B2(n17), .A(n29), .ZN(IMM[23]) );
  OAI21_X1 U47 ( .B1(n28), .B2(n16), .A(n29), .ZN(IMM[24]) );
  NOR2_X1 U48 ( .A1(n30), .A2(n42), .ZN(IMM[11]) );
  NOR2_X1 U49 ( .A1(n30), .A2(n41), .ZN(IMM[12]) );
  NOR2_X1 U50 ( .A1(n30), .A2(n40), .ZN(IMM[13]) );
  NOR2_X1 U51 ( .A1(n30), .A2(n39), .ZN(IMM[14]) );
  NOR2_X1 U52 ( .A1(n30), .A2(n38), .ZN(IMM[15]) );
  AND2_X1 U53 ( .A1(INST_IN[1]), .A2(n12), .ZN(IMM[1]) );
  AND2_X1 U55 ( .A1(INST_IN[3]), .A2(n12), .ZN(IMM[3]) );
  AND2_X1 U56 ( .A1(INST_IN[2]), .A2(n12), .ZN(IMM[2]) );
  AND2_X1 U57 ( .A1(INST_IN[5]), .A2(n12), .ZN(IMM[5]) );
  AND2_X1 U58 ( .A1(INST_IN[4]), .A2(n12), .ZN(IMM[4]) );
  AND2_X1 U59 ( .A1(INST_IN[6]), .A2(n12), .ZN(IMM[6]) );
  AND2_X1 U60 ( .A1(INST_IN[7]), .A2(n12), .ZN(IMM[7]) );
  AND2_X1 U61 ( .A1(INST_IN[8]), .A2(n12), .ZN(IMM[8]) );
  AND2_X1 U62 ( .A1(INST_IN[9]), .A2(n12), .ZN(IMM[9]) );
  AND2_X1 U63 ( .A1(INST_IN[10]), .A2(n12), .ZN(IMM[10]) );
  AND2_X1 U64 ( .A1(INST_IN[0]), .A2(n12), .ZN(IMM[0]) );
  INV_X1 U65 ( .A(INST_IN[23]), .ZN(n17) );
  INV_X1 U66 ( .A(n3), .ZN(RD2) );
  INV_X1 U67 ( .A(RD1), .ZN(n4) );
  AND2_X1 U68 ( .A1(n13), .A2(n35), .ZN(n6) );
  INV_X1 U69 ( .A(INST_IN[22]), .ZN(n18) );
  NOR2_X1 U70 ( .A1(n5), .A2(n23), .ZN(ADD_RS2[1]) );
  NOR2_X1 U71 ( .A1(n6), .A2(n21), .ZN(ADD_RS2[3]) );
  INV_X1 U72 ( .A(RD1), .ZN(n9) );
  INV_X1 U73 ( .A(INST_IN[24]), .ZN(n16) );
  NAND2_X1 U74 ( .A1(Jtype), .A2(n9), .ZN(n28) );
  NAND2_X1 U75 ( .A1(n1), .A2(n13), .ZN(n31) );
  OAI21_X1 U76 ( .B1(n1), .B2(Jtype), .A(n13), .ZN(n30) );
  INV_X1 U77 ( .A(INST_IN[29]), .ZN(n14) );
  NOR2_X1 U78 ( .A1(n10), .A2(n38), .ZN(n27) );
  AND3_X1 U79 ( .A1(Jtype), .A2(n10), .A3(INST_IN[25]), .ZN(n26) );
  INV_X1 U82 ( .A(n1), .ZN(n10) );
  INV_X1 U83 ( .A(INST_IN[27]), .ZN(n15) );
  NOR3_X1 U84 ( .A1(n14), .A2(INST_IN[30]), .A3(INST_IN[28]), .ZN(n37) );
  OR4_X1 U85 ( .A1(n15), .A2(INST_IN[28]), .A3(INST_IN[29]), .A4(INST_IN[31]), 
        .ZN(n33) );
  NAND4_X1 U86 ( .A1(Itype), .A2(INST_IN[31]), .A3(n36), .A4(n37), .ZN(n35) );
endmodule


module regn_N32_7 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U6 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U7 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U8 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U9 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U10 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U11 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U12 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U13 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U14 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U15 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U16 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U17 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U18 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U19 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U20 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U21 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U22 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U23 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U24 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U25 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U26 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U27 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U28 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U29 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U30 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U31 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U32 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U33 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U34 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U35 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U36 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U37 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U38 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U39 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U40 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U41 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U42 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U43 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U44 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U45 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U46 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U47 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U48 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U49 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U50 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U51 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U52 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U53 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U54 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U55 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U56 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U57 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U58 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U59 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U60 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U61 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U62 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U63 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U64 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U65 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U66 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module regn_N32_6 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U6 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U7 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U8 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U9 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U10 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U11 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U12 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U13 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U14 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U15 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U16 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U17 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U18 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  OAI21_X1 U19 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U20 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U21 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U22 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U23 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U24 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U25 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U26 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U27 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U28 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U29 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U30 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U31 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U32 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U33 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U34 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U35 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U36 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U37 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U38 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U39 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U40 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U41 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U42 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U43 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U44 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U45 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U46 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U47 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U48 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U49 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U50 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U51 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U52 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U53 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U54 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U55 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U56 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U57 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U58 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U59 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U60 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U61 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U62 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U63 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U64 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U65 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U66 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U67 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U68 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
endmodule


module regn_N5_0 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 DOUT_reg_4_ ( .D(n15), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n10) );
  DFFR_X1 DOUT_reg_3_ ( .D(n14), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n9) );
  DFFR_X1 DOUT_reg_2_ ( .D(n13), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n8) );
  DFFR_X1 DOUT_reg_1_ ( .D(n12), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n7) );
  DFFR_X1 DOUT_reg_0_ ( .D(n11), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n6) );
  OAI21_X1 U2 ( .B1(n7), .B2(EN), .A(n2), .ZN(n12) );
  NAND2_X1 U3 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U4 ( .B1(n8), .B2(EN), .A(n3), .ZN(n13) );
  NAND2_X1 U5 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U6 ( .B1(n9), .B2(EN), .A(n4), .ZN(n14) );
  NAND2_X1 U7 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U8 ( .B1(n10), .B2(EN), .A(n5), .ZN(n15) );
  NAND2_X1 U9 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U10 ( .B1(n6), .B2(EN), .A(n1), .ZN(n11) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
endmodule


module regn_N5_4 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 DOUT_reg_4_ ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21) );
  DFFR_X1 DOUT_reg_3_ ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22) );
  DFFR_X1 DOUT_reg_2_ ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23) );
  DFFR_X1 DOUT_reg_1_ ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24) );
  DFFR_X1 DOUT_reg_0_ ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U3 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
endmodule


module regn_N5_3 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 DOUT_reg_4_ ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21) );
  DFFR_X1 DOUT_reg_3_ ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22) );
  DFFR_X1 DOUT_reg_2_ ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23) );
  DFFR_X1 DOUT_reg_1_ ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24) );
  DFFR_X1 DOUT_reg_0_ ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U3 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
endmodule


module mux21_NBIT5_0 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n7, n8, n9, n10, n11, n1, n2, n3;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  INV_X1 U3 ( .A(n7), .ZN(Z[4]) );
  AOI22_X1 U4 ( .A1(A[4]), .A2(n3), .B1(n2), .B2(B[4]), .ZN(n7) );
  INV_X1 U5 ( .A(n10), .ZN(Z[1]) );
  INV_X1 U6 ( .A(n9), .ZN(Z[2]) );
  INV_X1 U7 ( .A(n8), .ZN(Z[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n1), .ZN(n8) );
  INV_X1 U9 ( .A(n11), .ZN(Z[0]) );
  AOI22_X1 U10 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n1), .ZN(n10) );
  AOI22_X1 U11 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n1), .ZN(n9) );
  AOI22_X1 U12 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n1), .ZN(n11) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module mux21_NBIT5_2 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n1, n2, n3, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  INV_X1 U3 ( .A(n18), .ZN(Z[4]) );
  INV_X1 U4 ( .A(n15), .ZN(Z[1]) );
  INV_X1 U5 ( .A(n16), .ZN(Z[2]) );
  INV_X1 U6 ( .A(n17), .ZN(Z[3]) );
  AOI22_X1 U7 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n1), .ZN(n17) );
  INV_X1 U8 ( .A(n14), .ZN(Z[0]) );
  AOI22_X1 U9 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n1), .ZN(n15) );
  AOI22_X1 U10 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n1), .ZN(n16) );
  AOI22_X1 U11 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n1), .ZN(n14) );
  AOI22_X1 U12 ( .A1(A[4]), .A2(n3), .B1(n2), .B2(B[4]), .ZN(n18) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module mux21_NBIT5_1 ( A, B, S, Z );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Z;
  input S;
  wire   n1, n2, n3, n14, n15, n16, n17, n18;

  BUF_X1 U1 ( .A(S), .Z(n1) );
  BUF_X1 U2 ( .A(S), .Z(n2) );
  INV_X1 U3 ( .A(n15), .ZN(Z[1]) );
  AOI22_X1 U4 ( .A1(A[1]), .A2(n3), .B1(B[1]), .B2(n1), .ZN(n15) );
  INV_X1 U5 ( .A(n16), .ZN(Z[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n3), .B1(B[2]), .B2(n1), .ZN(n16) );
  INV_X1 U7 ( .A(n17), .ZN(Z[3]) );
  AOI22_X1 U8 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(n1), .ZN(n17) );
  INV_X1 U9 ( .A(n18), .ZN(Z[4]) );
  AOI22_X1 U10 ( .A1(A[4]), .A2(n3), .B1(n2), .B2(B[4]), .ZN(n18) );
  INV_X1 U11 ( .A(n14), .ZN(Z[0]) );
  AOI22_X1 U12 ( .A1(A[0]), .A2(n3), .B1(B[0]), .B2(n1), .ZN(n14) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module register_file_NBIT_ADD5_NBIT_DATA32 ( CLK, RST, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RS1, ADD_RS2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, ENABLE, RD1, RD2, WR;
  wire   n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446;

  DFFR_X1 REGISTERS_reg_8__23_ ( .D(n3329), .CK(CLK), .RN(n665), .QN(n237) );
  DFFR_X1 REGISTERS_reg_8__22_ ( .D(n3328), .CK(CLK), .RN(n665), .QN(n238) );
  DFFR_X1 REGISTERS_reg_8__21_ ( .D(n3327), .CK(CLK), .RN(n665), .QN(n239) );
  DFFR_X1 REGISTERS_reg_8__20_ ( .D(n3326), .CK(CLK), .RN(n665), .QN(n240) );
  DFFR_X1 REGISTERS_reg_8__19_ ( .D(n3325), .CK(CLK), .RN(n665), .QN(n241) );
  DFFR_X1 REGISTERS_reg_8__18_ ( .D(n3324), .CK(CLK), .RN(n664), .QN(n242) );
  DFFR_X1 REGISTERS_reg_8__17_ ( .D(n3323), .CK(CLK), .RN(n664), .QN(n243) );
  DFFR_X1 REGISTERS_reg_8__16_ ( .D(n3322), .CK(CLK), .RN(n664), .QN(n244) );
  DFFR_X1 REGISTERS_reg_8__15_ ( .D(n3321), .CK(CLK), .RN(n664), .QN(n245) );
  DFFR_X1 REGISTERS_reg_8__14_ ( .D(n3320), .CK(CLK), .RN(n664), .QN(n246) );
  DFFR_X1 REGISTERS_reg_8__13_ ( .D(n3319), .CK(CLK), .RN(n664), .QN(n247) );
  DFFR_X1 REGISTERS_reg_8__12_ ( .D(n3318), .CK(CLK), .RN(n664), .QN(n248) );
  DFFR_X1 REGISTERS_reg_8__11_ ( .D(n3317), .CK(CLK), .RN(n664), .QN(n249) );
  DFFR_X1 REGISTERS_reg_8__10_ ( .D(n3316), .CK(CLK), .RN(n664), .QN(n250) );
  DFFR_X1 REGISTERS_reg_8__9_ ( .D(n3315), .CK(CLK), .RN(n664), .QN(n251) );
  DFFR_X1 REGISTERS_reg_8__8_ ( .D(n3314), .CK(CLK), .RN(n664), .QN(n252) );
  DFFR_X1 REGISTERS_reg_8__7_ ( .D(n3313), .CK(CLK), .RN(n669), .QN(n253) );
  DFFR_X1 REGISTERS_reg_8__6_ ( .D(n3312), .CK(CLK), .RN(n611), .QN(n254) );
  DFFR_X1 REGISTERS_reg_8__5_ ( .D(n3311), .CK(CLK), .RN(n611), .QN(n255) );
  DFFR_X1 REGISTERS_reg_8__4_ ( .D(n3310), .CK(CLK), .RN(n611), .QN(n256) );
  DFFR_X1 REGISTERS_reg_8__3_ ( .D(n3309), .CK(CLK), .RN(n611), .QN(n257) );
  DFFR_X1 REGISTERS_reg_8__2_ ( .D(n3308), .CK(CLK), .RN(n611), .QN(n258) );
  DFFR_X1 REGISTERS_reg_8__1_ ( .D(n3307), .CK(CLK), .RN(n610), .QN(n259) );
  DFFR_X1 REGISTERS_reg_8__0_ ( .D(n3306), .CK(CLK), .RN(n610), .QN(n260) );
  DFFR_X1 REGISTERS_reg_9__23_ ( .D(n3297), .CK(CLK), .RN(n610), .QN(n269) );
  DFFR_X1 REGISTERS_reg_9__22_ ( .D(n3296), .CK(CLK), .RN(n610), .QN(n270) );
  DFFR_X1 REGISTERS_reg_9__21_ ( .D(n3295), .CK(CLK), .RN(n609), .QN(n271) );
  DFFR_X1 REGISTERS_reg_9__20_ ( .D(n3294), .CK(CLK), .RN(n609), .QN(n272) );
  DFFR_X1 REGISTERS_reg_9__19_ ( .D(n3293), .CK(CLK), .RN(n609), .QN(n273) );
  DFFR_X1 REGISTERS_reg_9__18_ ( .D(n3292), .CK(CLK), .RN(n609), .QN(n274) );
  DFFR_X1 REGISTERS_reg_9__17_ ( .D(n3291), .CK(CLK), .RN(n609), .QN(n275) );
  DFFR_X1 REGISTERS_reg_9__16_ ( .D(n3290), .CK(CLK), .RN(n609), .QN(n276) );
  DFFR_X1 REGISTERS_reg_9__15_ ( .D(n3289), .CK(CLK), .RN(n609), .QN(n277) );
  DFFR_X1 REGISTERS_reg_9__14_ ( .D(n3288), .CK(CLK), .RN(n609), .QN(n278) );
  DFFR_X1 REGISTERS_reg_9__13_ ( .D(n3287), .CK(CLK), .RN(n609), .QN(n279) );
  DFFR_X1 REGISTERS_reg_9__12_ ( .D(n3286), .CK(CLK), .RN(n609), .QN(n280) );
  DFFR_X1 REGISTERS_reg_9__11_ ( .D(n3285), .CK(CLK), .RN(n609), .QN(n281) );
  DFFR_X1 REGISTERS_reg_9__10_ ( .D(n3284), .CK(CLK), .RN(n609), .QN(n282) );
  DFFR_X1 REGISTERS_reg_9__9_ ( .D(n3283), .CK(CLK), .RN(n608), .QN(n283) );
  DFFR_X1 REGISTERS_reg_9__8_ ( .D(n3282), .CK(CLK), .RN(n608), .QN(n284) );
  DFFR_X1 REGISTERS_reg_9__7_ ( .D(n3281), .CK(CLK), .RN(n608), .QN(n285) );
  DFFR_X1 REGISTERS_reg_9__6_ ( .D(n3280), .CK(CLK), .RN(n608), .QN(n286) );
  DFFR_X1 REGISTERS_reg_9__5_ ( .D(n3279), .CK(CLK), .RN(n608), .QN(n287) );
  DFFR_X1 REGISTERS_reg_9__4_ ( .D(n3278), .CK(CLK), .RN(n608), .QN(n288) );
  DFFR_X1 REGISTERS_reg_9__3_ ( .D(n3277), .CK(CLK), .RN(n608), .QN(n289) );
  DFFR_X1 REGISTERS_reg_9__2_ ( .D(n3276), .CK(CLK), .RN(n608), .QN(n290) );
  DFFR_X1 REGISTERS_reg_9__1_ ( .D(n3275), .CK(CLK), .RN(n608), .QN(n291) );
  DFFR_X1 REGISTERS_reg_9__0_ ( .D(n3274), .CK(CLK), .RN(n608), .QN(n292) );
  DFFR_X1 REGISTERS_reg_12__14_ ( .D(n3192), .CK(CLK), .RN(n601), .QN(n374) );
  DFFR_X1 REGISTERS_reg_12__13_ ( .D(n3191), .CK(CLK), .RN(n601), .QN(n375) );
  DFFR_X1 REGISTERS_reg_12__12_ ( .D(n3190), .CK(CLK), .RN(n601), .QN(n376) );
  DFFR_X1 REGISTERS_reg_12__11_ ( .D(n3189), .CK(CLK), .RN(n606), .QN(n377) );
  DFFR_X1 REGISTERS_reg_12__10_ ( .D(n3188), .CK(CLK), .RN(n653), .QN(n378) );
  DFFR_X1 REGISTERS_reg_12__9_ ( .D(n3187), .CK(CLK), .RN(n653), .QN(n379) );
  DFFR_X1 REGISTERS_reg_12__8_ ( .D(n3186), .CK(CLK), .RN(n653), .QN(n380) );
  DFFR_X1 REGISTERS_reg_12__7_ ( .D(n3185), .CK(CLK), .RN(n653), .QN(n381) );
  DFFR_X1 REGISTERS_reg_12__6_ ( .D(n3184), .CK(CLK), .RN(n653), .QN(n382) );
  DFFR_X1 REGISTERS_reg_12__5_ ( .D(n3183), .CK(CLK), .RN(n653), .QN(n383) );
  DFFR_X1 REGISTERS_reg_12__4_ ( .D(n3182), .CK(CLK), .RN(n653), .QN(n384) );
  DFFR_X1 REGISTERS_reg_12__3_ ( .D(n3181), .CK(CLK), .RN(n653), .QN(n385) );
  DFFR_X1 REGISTERS_reg_12__2_ ( .D(n3180), .CK(CLK), .RN(n652), .QN(n386) );
  DFFR_X1 REGISTERS_reg_12__1_ ( .D(n3179), .CK(CLK), .RN(n652), .QN(n387) );
  DFFR_X1 REGISTERS_reg_12__0_ ( .D(n3178), .CK(CLK), .RN(n652), .QN(n388) );
  DFFR_X1 REGISTERS_reg_17__23_ ( .D(n3041), .CK(CLK), .RN(n703), .QN(n525) );
  DFFR_X1 REGISTERS_reg_17__22_ ( .D(n3040), .CK(CLK), .RN(n703), .QN(n526) );
  DFFR_X1 REGISTERS_reg_17__21_ ( .D(n3039), .CK(CLK), .RN(n703), .QN(n527) );
  DFFR_X1 REGISTERS_reg_17__20_ ( .D(n3038), .CK(CLK), .RN(n703), .QN(n528) );
  DFFR_X1 REGISTERS_reg_17__19_ ( .D(n3037), .CK(CLK), .RN(n703), .QN(n529) );
  DFFR_X1 REGISTERS_reg_17__18_ ( .D(n3036), .CK(CLK), .RN(n703), .QN(n530) );
  DFFR_X1 REGISTERS_reg_17__17_ ( .D(n3035), .CK(CLK), .RN(n702), .QN(n531) );
  DFFR_X1 REGISTERS_reg_17__16_ ( .D(n3034), .CK(CLK), .RN(n702), .QN(n532) );
  DFFR_X1 REGISTERS_reg_17__15_ ( .D(n3033), .CK(CLK), .RN(n702), .QN(n533) );
  DFFR_X1 REGISTERS_reg_17__14_ ( .D(n3032), .CK(CLK), .RN(n702), .QN(n534) );
  DFFR_X1 REGISTERS_reg_17__13_ ( .D(n3031), .CK(CLK), .RN(n702), .QN(n535) );
  DFFR_X1 REGISTERS_reg_17__12_ ( .D(n3030), .CK(CLK), .RN(n702), .QN(n536) );
  DFFR_X1 REGISTERS_reg_17__11_ ( .D(n3029), .CK(CLK), .RN(n702), .QN(n537) );
  DFFR_X1 REGISTERS_reg_17__10_ ( .D(n3028), .CK(CLK), .RN(n702), .QN(n538) );
  DFFR_X1 REGISTERS_reg_17__9_ ( .D(n3027), .CK(CLK), .RN(n702), .QN(n539) );
  DFFR_X1 REGISTERS_reg_17__8_ ( .D(n3026), .CK(CLK), .RN(n702), .QN(n540) );
  DFFR_X1 REGISTERS_reg_17__7_ ( .D(n3025), .CK(CLK), .RN(n702), .QN(n541) );
  DFFR_X1 REGISTERS_reg_17__6_ ( .D(n3024), .CK(CLK), .RN(n702), .QN(n542) );
  DFFR_X1 REGISTERS_reg_17__5_ ( .D(n3023), .CK(CLK), .RN(n701), .QN(n543) );
  DFFR_X1 REGISTERS_reg_17__4_ ( .D(n3022), .CK(CLK), .RN(n701), .QN(n544) );
  DFFR_X1 REGISTERS_reg_17__3_ ( .D(n3021), .CK(CLK), .RN(n701), .QN(n545) );
  DFFR_X1 REGISTERS_reg_17__2_ ( .D(n3020), .CK(CLK), .RN(n701), .QN(n546) );
  DFFR_X1 REGISTERS_reg_17__1_ ( .D(n3019), .CK(CLK), .RN(n701), .QN(n547) );
  DFFR_X1 REGISTERS_reg_17__0_ ( .D(n3018), .CK(CLK), .RN(n701), .QN(n548) );
  DFFR_X1 REGISTERS_reg_20__23_ ( .D(n2945), .CK(CLK), .RN(n695), .QN(n621) );
  DFFR_X1 REGISTERS_reg_20__22_ ( .D(n2944), .CK(CLK), .RN(n695), .QN(n622) );
  DFFR_X1 REGISTERS_reg_20__21_ ( .D(n2943), .CK(CLK), .RN(n695), .QN(n623) );
  DFFR_X1 REGISTERS_reg_20__20_ ( .D(n2942), .CK(CLK), .RN(n695), .QN(n624) );
  DFFR_X1 REGISTERS_reg_20__19_ ( .D(n2941), .CK(CLK), .RN(n700), .QN(n625) );
  DFFR_X1 REGISTERS_reg_20__18_ ( .D(n2940), .CK(CLK), .RN(n715), .QN(n626) );
  DFFR_X1 REGISTERS_reg_20__17_ ( .D(n2939), .CK(CLK), .RN(n715), .QN(n627) );
  DFFR_X1 REGISTERS_reg_20__16_ ( .D(n2938), .CK(CLK), .RN(n715), .QN(n628) );
  DFFR_X1 REGISTERS_reg_20__15_ ( .D(n2937), .CK(CLK), .RN(n715), .QN(n629) );
  DFFR_X1 REGISTERS_reg_20__14_ ( .D(n2936), .CK(CLK), .RN(n715), .QN(n630) );
  DFFR_X1 REGISTERS_reg_20__13_ ( .D(n2935), .CK(CLK), .RN(n715), .QN(n631) );
  DFFR_X1 REGISTERS_reg_20__12_ ( .D(n2934), .CK(CLK), .RN(n715), .QN(n632) );
  DFFR_X1 REGISTERS_reg_20__11_ ( .D(n2933), .CK(CLK), .RN(n715), .QN(n633) );
  DFFR_X1 REGISTERS_reg_20__10_ ( .D(n2932), .CK(CLK), .RN(n714), .QN(n634) );
  DFFR_X1 REGISTERS_reg_20__9_ ( .D(n2931), .CK(CLK), .RN(n714), .QN(n635) );
  DFFR_X1 REGISTERS_reg_20__8_ ( .D(n2930), .CK(CLK), .RN(n714), .QN(n636) );
  DFFR_X1 REGISTERS_reg_20__7_ ( .D(n2929), .CK(CLK), .RN(n714), .QN(n637) );
  DFFR_X1 REGISTERS_reg_20__6_ ( .D(n2928), .CK(CLK), .RN(n714), .QN(n638) );
  DFFR_X1 REGISTERS_reg_20__5_ ( .D(n2927), .CK(CLK), .RN(n714), .QN(n639) );
  DFFR_X1 REGISTERS_reg_20__4_ ( .D(n2926), .CK(CLK), .RN(n714), .QN(n640) );
  DFFR_X1 REGISTERS_reg_20__3_ ( .D(n2925), .CK(CLK), .RN(n714), .QN(n641) );
  DFFR_X1 REGISTERS_reg_20__2_ ( .D(n2924), .CK(CLK), .RN(n714), .QN(n642) );
  DFFR_X1 REGISTERS_reg_20__1_ ( .D(n2923), .CK(CLK), .RN(n714), .QN(n643) );
  DFFR_X1 REGISTERS_reg_20__0_ ( .D(n2922), .CK(CLK), .RN(n714), .QN(n644) );
  DFFR_X1 REGISTERS_reg_24__3_ ( .D(n2797), .CK(CLK), .RN(n683), .Q(n4034) );
  DFFR_X1 REGISTERS_reg_24__2_ ( .D(n2796), .CK(CLK), .RN(n682), .Q(n4033) );
  DFFR_X1 REGISTERS_reg_24__1_ ( .D(n2795), .CK(CLK), .RN(n682), .Q(n4032) );
  DFFR_X1 REGISTERS_reg_24__0_ ( .D(n2794), .CK(CLK), .RN(n682), .Q(n4031) );
  DFFR_X1 REGISTERS_reg_27__23_ ( .D(n2721), .CK(CLK), .RN(n676), .QN(n845) );
  DFFR_X1 REGISTERS_reg_27__22_ ( .D(n2720), .CK(CLK), .RN(n676), .QN(n846) );
  DFFR_X1 REGISTERS_reg_27__21_ ( .D(n2719), .CK(CLK), .RN(n676), .QN(n847) );
  DFFR_X1 REGISTERS_reg_27__20_ ( .D(n2718), .CK(CLK), .RN(n676), .QN(n848) );
  DFFR_X1 REGISTERS_reg_27__19_ ( .D(n2717), .CK(CLK), .RN(n676), .QN(n849) );
  DFFR_X1 REGISTERS_reg_27__18_ ( .D(n2716), .CK(CLK), .RN(n676), .QN(n850) );
  DFFR_X1 REGISTERS_reg_27__17_ ( .D(n2715), .CK(CLK), .RN(n676), .QN(n851) );
  DFFR_X1 REGISTERS_reg_27__16_ ( .D(n2714), .CK(CLK), .RN(n676), .QN(n852) );
  DFFR_X1 REGISTERS_reg_27__15_ ( .D(n2713), .CK(CLK), .RN(n675), .QN(n853) );
  DFFR_X1 REGISTERS_reg_27__14_ ( .D(n2712), .CK(CLK), .RN(n675), .QN(n854) );
  DFFR_X1 REGISTERS_reg_27__13_ ( .D(n2711), .CK(CLK), .RN(n675), .QN(n855) );
  DFFR_X1 REGISTERS_reg_27__12_ ( .D(n2710), .CK(CLK), .RN(n675), .QN(n856) );
  DFFR_X1 REGISTERS_reg_27__11_ ( .D(n2709), .CK(CLK), .RN(n675), .QN(n857) );
  DFFR_X1 REGISTERS_reg_27__10_ ( .D(n2708), .CK(CLK), .RN(n675), .QN(n858) );
  DFFR_X1 REGISTERS_reg_27__9_ ( .D(n2707), .CK(CLK), .RN(n675), .QN(n859) );
  DFFR_X1 REGISTERS_reg_27__8_ ( .D(n2706), .CK(CLK), .RN(n675), .QN(n860) );
  DFFR_X1 REGISTERS_reg_27__7_ ( .D(n2705), .CK(CLK), .RN(n675), .QN(n861) );
  DFFR_X1 REGISTERS_reg_27__6_ ( .D(n2704), .CK(CLK), .RN(n675), .QN(n862) );
  DFFR_X1 REGISTERS_reg_27__5_ ( .D(n2703), .CK(CLK), .RN(n675), .QN(n863) );
  DFFR_X1 REGISTERS_reg_27__4_ ( .D(n2702), .CK(CLK), .RN(n675), .QN(n864) );
  DFFR_X1 REGISTERS_reg_27__3_ ( .D(n2701), .CK(CLK), .RN(n674), .QN(n865) );
  DFFR_X1 REGISTERS_reg_27__2_ ( .D(n2700), .CK(CLK), .RN(n674), .QN(n866) );
  DFFR_X1 REGISTERS_reg_27__1_ ( .D(n2699), .CK(CLK), .RN(n674), .QN(n867) );
  DFFR_X1 REGISTERS_reg_27__0_ ( .D(n2698), .CK(CLK), .RN(n674), .QN(n868) );
  DFFR_X1 REGISTERS_reg_30__23_ ( .D(n2625), .CK(CLK), .RN(n689), .QN(n941) );
  DFFR_X1 REGISTERS_reg_30__22_ ( .D(n2624), .CK(CLK), .RN(n689), .QN(n942) );
  DFFR_X1 REGISTERS_reg_30__21_ ( .D(n2623), .CK(CLK), .RN(n689), .QN(n943) );
  DFFR_X1 REGISTERS_reg_30__20_ ( .D(n2622), .CK(CLK), .RN(n689), .QN(n944) );
  DFFR_X1 REGISTERS_reg_30__19_ ( .D(n2621), .CK(CLK), .RN(n688), .QN(n945) );
  DFFR_X1 REGISTERS_reg_30__18_ ( .D(n2620), .CK(CLK), .RN(n688), .QN(n946) );
  DFFR_X1 REGISTERS_reg_30__17_ ( .D(n2619), .CK(CLK), .RN(n688), .QN(n947) );
  DFFR_X1 REGISTERS_reg_30__16_ ( .D(n2618), .CK(CLK), .RN(n688), .QN(n948) );
  DFFR_X1 REGISTERS_reg_30__15_ ( .D(n2617), .CK(CLK), .RN(n688), .QN(n949) );
  DFFR_X1 REGISTERS_reg_30__14_ ( .D(n2616), .CK(CLK), .RN(n688), .QN(n950) );
  DFFR_X1 REGISTERS_reg_30__13_ ( .D(n2615), .CK(CLK), .RN(n688), .QN(n951) );
  DFFR_X1 REGISTERS_reg_30__12_ ( .D(n2614), .CK(CLK), .RN(n688), .QN(n952) );
  DFFR_X1 REGISTERS_reg_30__11_ ( .D(n2613), .CK(CLK), .RN(n688), .QN(n953) );
  DFFR_X1 REGISTERS_reg_30__10_ ( .D(n2612), .CK(CLK), .RN(n688), .QN(n954) );
  DFFR_X1 REGISTERS_reg_30__9_ ( .D(n2611), .CK(CLK), .RN(n688), .QN(n955) );
  DFFR_X1 REGISTERS_reg_30__8_ ( .D(n2610), .CK(CLK), .RN(n688), .QN(n956) );
  DFFR_X1 REGISTERS_reg_30__7_ ( .D(n2609), .CK(CLK), .RN(n687), .QN(n957) );
  DFFR_X1 REGISTERS_reg_30__6_ ( .D(n2608), .CK(CLK), .RN(n687), .QN(n958) );
  DFFR_X1 REGISTERS_reg_30__5_ ( .D(n2607), .CK(CLK), .RN(n687), .QN(n959) );
  DFFR_X1 REGISTERS_reg_30__4_ ( .D(n2606), .CK(CLK), .RN(n687), .QN(n960) );
  DFFR_X1 REGISTERS_reg_30__3_ ( .D(n2605), .CK(CLK), .RN(n687), .QN(n961) );
  DFFR_X1 REGISTERS_reg_30__2_ ( .D(n2604), .CK(CLK), .RN(n687), .QN(n962) );
  DFFR_X1 REGISTERS_reg_30__1_ ( .D(n2603), .CK(CLK), .RN(n687), .QN(n963) );
  DFFR_X1 REGISTERS_reg_30__0_ ( .D(n2602), .CK(CLK), .RN(n687), .QN(n964) );
  DFFR_X1 REGISTERS_reg_5__31_ ( .D(n3433), .CK(CLK), .RN(RST), .Q(n803) );
  DFFR_X1 REGISTERS_reg_5__30_ ( .D(n3432), .CK(CLK), .RN(n674), .Q(n805) );
  DFFR_X1 REGISTERS_reg_5__29_ ( .D(n3431), .CK(CLK), .RN(n673), .Q(n806) );
  DFFR_X1 REGISTERS_reg_5__28_ ( .D(n3430), .CK(CLK), .RN(n673), .Q(n807) );
  DFFR_X1 REGISTERS_reg_5__27_ ( .D(n3429), .CK(CLK), .RN(n673), .Q(n808) );
  DFFR_X1 REGISTERS_reg_5__26_ ( .D(n3428), .CK(CLK), .RN(n673), .Q(n809) );
  DFFR_X1 REGISTERS_reg_5__25_ ( .D(n3427), .CK(CLK), .RN(n673), .Q(n810) );
  DFFR_X1 REGISTERS_reg_5__24_ ( .D(n3426), .CK(CLK), .RN(n673), .Q(n811) );
  DFFR_X1 REGISTERS_reg_4__31_ ( .D(n3465), .CK(CLK), .RN(n656), .Q(n769) );
  DFFR_X1 REGISTERS_reg_4__30_ ( .D(n3464), .CK(CLK), .RN(n656), .Q(n771) );
  DFFR_X1 REGISTERS_reg_4__29_ ( .D(n3463), .CK(CLK), .RN(n655), .Q(n772) );
  DFFR_X1 REGISTERS_reg_4__28_ ( .D(n3462), .CK(CLK), .RN(n655), .Q(n773) );
  DFFR_X1 REGISTERS_reg_4__27_ ( .D(n3461), .CK(CLK), .RN(n655), .Q(n774) );
  DFFR_X1 REGISTERS_reg_4__26_ ( .D(n3460), .CK(CLK), .RN(n655), .Q(n775) );
  DFFR_X1 REGISTERS_reg_4__25_ ( .D(n3459), .CK(CLK), .RN(n655), .Q(n776) );
  DFFR_X1 REGISTERS_reg_4__24_ ( .D(n3458), .CK(CLK), .RN(n655), .Q(n777) );
  DFFR_X1 REGISTERS_reg_1__31_ ( .D(n3561), .CK(CLK), .RN(n674), .Q(n730) );
  DFFR_X1 REGISTERS_reg_1__30_ ( .D(n3560), .CK(CLK), .RN(n601), .Q(n732) );
  DFFR_X1 REGISTERS_reg_1__29_ ( .D(n3559), .CK(CLK), .RN(n664), .Q(n733) );
  DFFR_X1 REGISTERS_reg_1__28_ ( .D(n3558), .CK(CLK), .RN(n663), .Q(n734) );
  DFFR_X1 REGISTERS_reg_1__27_ ( .D(n3557), .CK(CLK), .RN(n663), .Q(n735) );
  DFFR_X1 REGISTERS_reg_1__26_ ( .D(n3556), .CK(CLK), .RN(n663), .Q(n736) );
  DFFR_X1 REGISTERS_reg_1__25_ ( .D(n3555), .CK(CLK), .RN(n663), .Q(n737) );
  DFFR_X1 REGISTERS_reg_1__24_ ( .D(n3554), .CK(CLK), .RN(n663), .Q(n738) );
  DFFR_X1 REGISTERS_reg_21__31_ ( .D(n2921), .CK(CLK), .RN(n714), .Q(n1148) );
  DFFR_X1 REGISTERS_reg_21__30_ ( .D(n2920), .CK(CLK), .RN(n713), .Q(n1150) );
  DFFR_X1 REGISTERS_reg_21__29_ ( .D(n2919), .CK(CLK), .RN(n713), .Q(n1151) );
  DFFR_X1 REGISTERS_reg_21__28_ ( .D(n2918), .CK(CLK), .RN(n713), .Q(n1152) );
  DFFR_X1 REGISTERS_reg_21__27_ ( .D(n2917), .CK(CLK), .RN(n713), .Q(n1153) );
  DFFR_X1 REGISTERS_reg_21__26_ ( .D(n2916), .CK(CLK), .RN(n713), .Q(n1154) );
  DFFR_X1 REGISTERS_reg_21__25_ ( .D(n2915), .CK(CLK), .RN(n713), .Q(n1155) );
  DFFR_X1 REGISTERS_reg_21__24_ ( .D(n2914), .CK(CLK), .RN(n713), .Q(n1156) );
  DFFR_X1 REGISTERS_reg_16__31_ ( .D(n3081), .CK(CLK), .RN(n612), .Q(n1046) );
  DFFR_X1 REGISTERS_reg_16__30_ ( .D(n3080), .CK(CLK), .RN(n612), .Q(n1048) );
  DFFR_X1 REGISTERS_reg_16__29_ ( .D(n3079), .CK(CLK), .RN(n612), .Q(n1049) );
  DFFR_X1 REGISTERS_reg_16__28_ ( .D(n3078), .CK(CLK), .RN(n612), .Q(n1050) );
  DFFR_X1 REGISTERS_reg_16__27_ ( .D(n3077), .CK(CLK), .RN(n612), .Q(n1051) );
  DFFR_X1 REGISTERS_reg_16__26_ ( .D(n3076), .CK(CLK), .RN(n612), .Q(n1052) );
  DFFR_X1 REGISTERS_reg_16__25_ ( .D(n3075), .CK(CLK), .RN(n612), .Q(n1053) );
  DFFR_X1 REGISTERS_reg_16__24_ ( .D(n3074), .CK(CLK), .RN(n612), .Q(n1054) );
  DFFR_X1 REGISTERS_reg_31__31_ ( .D(n2601), .CK(CLK), .RN(n687), .Q(n1289) );
  DFFR_X1 REGISTERS_reg_31__30_ ( .D(n2600), .CK(CLK), .RN(n687), .Q(n1291) );
  DFFR_X1 REGISTERS_reg_31__29_ ( .D(n2599), .CK(CLK), .RN(n687), .Q(n1292) );
  DFFR_X1 REGISTERS_reg_31__28_ ( .D(n2598), .CK(CLK), .RN(n687), .Q(n1293) );
  DFFR_X1 REGISTERS_reg_31__27_ ( .D(n2597), .CK(CLK), .RN(n686), .Q(n1294) );
  DFFR_X1 REGISTERS_reg_31__26_ ( .D(n2596), .CK(CLK), .RN(n686), .Q(n1295) );
  DFFR_X1 REGISTERS_reg_31__25_ ( .D(n2595), .CK(CLK), .RN(n686), .Q(n1296) );
  DFFR_X1 REGISTERS_reg_31__24_ ( .D(n2594), .CK(CLK), .RN(n686), .Q(n1297) );
  DFFR_X1 REGISTERS_reg_26__31_ ( .D(n2761), .CK(CLK), .RN(n680), .Q(n1187) );
  DFFR_X1 REGISTERS_reg_26__30_ ( .D(n2760), .CK(CLK), .RN(n679), .Q(n1189) );
  DFFR_X1 REGISTERS_reg_26__29_ ( .D(n2759), .CK(CLK), .RN(n679), .Q(n1190) );
  DFFR_X1 REGISTERS_reg_26__28_ ( .D(n2758), .CK(CLK), .RN(n679), .Q(n1191) );
  DFFR_X1 REGISTERS_reg_26__27_ ( .D(n2757), .CK(CLK), .RN(n679), .Q(n1192) );
  DFFR_X1 REGISTERS_reg_26__26_ ( .D(n2756), .CK(CLK), .RN(n679), .Q(n1193) );
  DFFR_X1 REGISTERS_reg_26__25_ ( .D(n2755), .CK(CLK), .RN(n679), .Q(n1194) );
  DFFR_X1 REGISTERS_reg_26__24_ ( .D(n2754), .CK(CLK), .RN(n679), .Q(n1195) );
  DFFR_X1 REGISTERS_reg_5__23_ ( .D(n3425), .CK(CLK), .RN(n673), .Q(n812) );
  DFFR_X1 REGISTERS_reg_5__22_ ( .D(n3424), .CK(CLK), .RN(n673), .Q(n813) );
  DFFR_X1 REGISTERS_reg_5__21_ ( .D(n3423), .CK(CLK), .RN(n673), .Q(n814) );
  DFFR_X1 REGISTERS_reg_5__20_ ( .D(n3422), .CK(CLK), .RN(n673), .Q(n815) );
  DFFR_X1 REGISTERS_reg_5__19_ ( .D(n3421), .CK(CLK), .RN(n673), .Q(n816) );
  DFFR_X1 REGISTERS_reg_5__18_ ( .D(n3420), .CK(CLK), .RN(n673), .Q(n817) );
  DFFR_X1 REGISTERS_reg_5__17_ ( .D(n3419), .CK(CLK), .RN(n672), .Q(n818) );
  DFFR_X1 REGISTERS_reg_5__16_ ( .D(n3418), .CK(CLK), .RN(n672), .Q(n819) );
  DFFR_X1 REGISTERS_reg_5__15_ ( .D(n3417), .CK(CLK), .RN(n672), .Q(n820) );
  DFFR_X1 REGISTERS_reg_5__14_ ( .D(n3416), .CK(CLK), .RN(n672), .Q(n821) );
  DFFR_X1 REGISTERS_reg_5__13_ ( .D(n3415), .CK(CLK), .RN(n672), .Q(n822) );
  DFFR_X1 REGISTERS_reg_5__12_ ( .D(n3414), .CK(CLK), .RN(n672), .Q(n823) );
  DFFR_X1 REGISTERS_reg_5__11_ ( .D(n3413), .CK(CLK), .RN(n672), .Q(n824) );
  DFFR_X1 REGISTERS_reg_5__10_ ( .D(n3412), .CK(CLK), .RN(n672), .Q(n825) );
  DFFR_X1 REGISTERS_reg_5__9_ ( .D(n3411), .CK(CLK), .RN(n672), .Q(n826) );
  DFFR_X1 REGISTERS_reg_5__8_ ( .D(n3410), .CK(CLK), .RN(n672), .Q(n827) );
  DFFR_X1 REGISTERS_reg_5__7_ ( .D(n3409), .CK(CLK), .RN(n672), .Q(n828) );
  DFFR_X1 REGISTERS_reg_5__6_ ( .D(n3408), .CK(CLK), .RN(n672), .Q(n829) );
  DFFR_X1 REGISTERS_reg_5__5_ ( .D(n3407), .CK(CLK), .RN(n671), .Q(n830) );
  DFFR_X1 REGISTERS_reg_5__4_ ( .D(n3406), .CK(CLK), .RN(n671), .Q(n831) );
  DFFR_X1 REGISTERS_reg_5__3_ ( .D(n3405), .CK(CLK), .RN(n671), .Q(n832) );
  DFFR_X1 REGISTERS_reg_5__2_ ( .D(n3404), .CK(CLK), .RN(n671), .Q(n833) );
  DFFR_X1 REGISTERS_reg_5__1_ ( .D(n3403), .CK(CLK), .RN(n671), .Q(n834) );
  DFFR_X1 REGISTERS_reg_5__0_ ( .D(n3402), .CK(CLK), .RN(n671), .Q(n835) );
  DFFR_X1 REGISTERS_reg_4__23_ ( .D(n3457), .CK(CLK), .RN(n655), .Q(n778) );
  DFFR_X1 REGISTERS_reg_4__22_ ( .D(n3456), .CK(CLK), .RN(n655), .Q(n779) );
  DFFR_X1 REGISTERS_reg_4__21_ ( .D(n3455), .CK(CLK), .RN(n655), .Q(n780) );
  DFFR_X1 REGISTERS_reg_4__20_ ( .D(n3454), .CK(CLK), .RN(n655), .Q(n781) );
  DFFR_X1 REGISTERS_reg_4__19_ ( .D(n3453), .CK(CLK), .RN(n655), .Q(n782) );
  DFFR_X1 REGISTERS_reg_4__18_ ( .D(n3452), .CK(CLK), .RN(n655), .Q(n783) );
  DFFR_X1 REGISTERS_reg_4__17_ ( .D(n3451), .CK(CLK), .RN(n654), .Q(n784) );
  DFFR_X1 REGISTERS_reg_4__16_ ( .D(n3450), .CK(CLK), .RN(n654), .Q(n785) );
  DFFR_X1 REGISTERS_reg_4__15_ ( .D(n3449), .CK(CLK), .RN(n654), .Q(n786) );
  DFFR_X1 REGISTERS_reg_4__14_ ( .D(n3448), .CK(CLK), .RN(n654), .Q(n787) );
  DFFR_X1 REGISTERS_reg_4__13_ ( .D(n3447), .CK(CLK), .RN(n654), .Q(n788) );
  DFFR_X1 REGISTERS_reg_4__12_ ( .D(n3446), .CK(CLK), .RN(n654), .Q(n789) );
  DFFR_X1 REGISTERS_reg_4__11_ ( .D(n3445), .CK(CLK), .RN(n654), .Q(n790) );
  DFFR_X1 REGISTERS_reg_4__10_ ( .D(n3444), .CK(CLK), .RN(n654), .Q(n791) );
  DFFR_X1 REGISTERS_reg_4__9_ ( .D(n3443), .CK(CLK), .RN(n654), .Q(n792) );
  DFFR_X1 REGISTERS_reg_4__8_ ( .D(n3442), .CK(CLK), .RN(n654), .Q(n793) );
  DFFR_X1 REGISTERS_reg_4__7_ ( .D(n3441), .CK(CLK), .RN(n654), .Q(n794) );
  DFFR_X1 REGISTERS_reg_4__6_ ( .D(n3440), .CK(CLK), .RN(n654), .Q(n795) );
  DFFR_X1 REGISTERS_reg_4__5_ ( .D(n3439), .CK(CLK), .RN(n653), .Q(n796) );
  DFFR_X1 REGISTERS_reg_4__4_ ( .D(n3438), .CK(CLK), .RN(n653), .Q(n797) );
  DFFR_X1 REGISTERS_reg_4__3_ ( .D(n3437), .CK(CLK), .RN(n653), .Q(n798) );
  DFFR_X1 REGISTERS_reg_4__2_ ( .D(n3436), .CK(CLK), .RN(n658), .Q(n799) );
  DFFR_X1 REGISTERS_reg_4__1_ ( .D(n3435), .CK(CLK), .RN(n674), .Q(n800) );
  DFFR_X1 REGISTERS_reg_4__0_ ( .D(n3434), .CK(CLK), .RN(n674), .Q(n801) );
  DFFR_X1 REGISTERS_reg_1__23_ ( .D(n3553), .CK(CLK), .RN(n663), .Q(n739) );
  DFFR_X1 REGISTERS_reg_1__22_ ( .D(n3552), .CK(CLK), .RN(n663), .Q(n740) );
  DFFR_X1 REGISTERS_reg_1__21_ ( .D(n3551), .CK(CLK), .RN(n663), .Q(n741) );
  DFFR_X1 REGISTERS_reg_1__20_ ( .D(n3550), .CK(CLK), .RN(n663), .Q(n742) );
  DFFR_X1 REGISTERS_reg_1__19_ ( .D(n3549), .CK(CLK), .RN(n663), .Q(n743) );
  DFFR_X1 REGISTERS_reg_1__18_ ( .D(n3548), .CK(CLK), .RN(n663), .Q(n744) );
  DFFR_X1 REGISTERS_reg_1__17_ ( .D(n3547), .CK(CLK), .RN(n663), .Q(n745) );
  DFFR_X1 REGISTERS_reg_1__16_ ( .D(n3546), .CK(CLK), .RN(n662), .Q(n746) );
  DFFR_X1 REGISTERS_reg_1__15_ ( .D(n3545), .CK(CLK), .RN(n662), .Q(n747) );
  DFFR_X1 REGISTERS_reg_1__14_ ( .D(n3544), .CK(CLK), .RN(n662), .Q(n748) );
  DFFR_X1 REGISTERS_reg_1__13_ ( .D(n3543), .CK(CLK), .RN(n662), .Q(n749) );
  DFFR_X1 REGISTERS_reg_1__12_ ( .D(n3542), .CK(CLK), .RN(n662), .Q(n750) );
  DFFR_X1 REGISTERS_reg_1__11_ ( .D(n3541), .CK(CLK), .RN(n662), .Q(n751) );
  DFFR_X1 REGISTERS_reg_1__10_ ( .D(n3540), .CK(CLK), .RN(n662), .Q(n752) );
  DFFR_X1 REGISTERS_reg_1__9_ ( .D(n3539), .CK(CLK), .RN(n662), .Q(n753) );
  DFFR_X1 REGISTERS_reg_1__8_ ( .D(n3538), .CK(CLK), .RN(n662), .Q(n754) );
  DFFR_X1 REGISTERS_reg_1__7_ ( .D(n3537), .CK(CLK), .RN(n662), .Q(n755) );
  DFFR_X1 REGISTERS_reg_1__6_ ( .D(n3536), .CK(CLK), .RN(n662), .Q(n756) );
  DFFR_X1 REGISTERS_reg_1__5_ ( .D(n3535), .CK(CLK), .RN(n662), .Q(n757) );
  DFFR_X1 REGISTERS_reg_1__4_ ( .D(n3534), .CK(CLK), .RN(n661), .Q(n758) );
  DFFR_X1 REGISTERS_reg_1__3_ ( .D(n3533), .CK(CLK), .RN(n661), .Q(n759) );
  DFFR_X1 REGISTERS_reg_1__2_ ( .D(n3532), .CK(CLK), .RN(n661), .Q(n760) );
  DFFR_X1 REGISTERS_reg_1__1_ ( .D(n3531), .CK(CLK), .RN(n661), .Q(n761) );
  DFFR_X1 REGISTERS_reg_1__0_ ( .D(n3530), .CK(CLK), .RN(n661), .Q(n762) );
  DFFR_X1 REGISTERS_reg_13__31_ ( .D(n3177), .CK(CLK), .RN(n652), .QN(n389) );
  DFFR_X1 REGISTERS_reg_13__30_ ( .D(n3176), .CK(CLK), .RN(n652), .QN(n390) );
  DFFR_X1 REGISTERS_reg_13__29_ ( .D(n3175), .CK(CLK), .RN(n652), .QN(n391) );
  DFFR_X1 REGISTERS_reg_13__28_ ( .D(n3174), .CK(CLK), .RN(n652), .QN(n392) );
  DFFR_X1 REGISTERS_reg_13__27_ ( .D(n3173), .CK(CLK), .RN(n652), .QN(n393) );
  DFFR_X1 REGISTERS_reg_13__26_ ( .D(n3172), .CK(CLK), .RN(n652), .QN(n394) );
  DFFR_X1 REGISTERS_reg_13__25_ ( .D(n3171), .CK(CLK), .RN(n652), .QN(n395) );
  DFFR_X1 REGISTERS_reg_13__24_ ( .D(n3170), .CK(CLK), .RN(n652), .QN(n396) );
  DFFR_X1 REGISTERS_reg_12__31_ ( .D(n3209), .CK(CLK), .RN(n602), .QN(n357) );
  DFFR_X1 REGISTERS_reg_12__30_ ( .D(n3208), .CK(CLK), .RN(n602), .QN(n358) );
  DFFR_X1 REGISTERS_reg_12__29_ ( .D(n3207), .CK(CLK), .RN(n602), .QN(n359) );
  DFFR_X1 REGISTERS_reg_12__28_ ( .D(n3206), .CK(CLK), .RN(n602), .QN(n360) );
  DFFR_X1 REGISTERS_reg_12__27_ ( .D(n3205), .CK(CLK), .RN(n602), .QN(n361) );
  DFFR_X1 REGISTERS_reg_12__26_ ( .D(n3204), .CK(CLK), .RN(n602), .QN(n362) );
  DFFR_X1 REGISTERS_reg_12__25_ ( .D(n3203), .CK(CLK), .RN(n602), .QN(n363) );
  DFFR_X1 REGISTERS_reg_12__24_ ( .D(n3202), .CK(CLK), .RN(n602), .QN(n364) );
  DFFR_X1 REGISTERS_reg_20__31_ ( .D(n2953), .CK(CLK), .RN(n696), .QN(n613) );
  DFFR_X1 REGISTERS_reg_20__30_ ( .D(n2952), .CK(CLK), .RN(n695), .QN(n614) );
  DFFR_X1 REGISTERS_reg_20__29_ ( .D(n2951), .CK(CLK), .RN(n695), .QN(n615) );
  DFFR_X1 REGISTERS_reg_20__28_ ( .D(n2950), .CK(CLK), .RN(n695), .QN(n616) );
  DFFR_X1 REGISTERS_reg_20__27_ ( .D(n2949), .CK(CLK), .RN(n695), .QN(n617) );
  DFFR_X1 REGISTERS_reg_20__26_ ( .D(n2948), .CK(CLK), .RN(n695), .QN(n618) );
  DFFR_X1 REGISTERS_reg_20__25_ ( .D(n2947), .CK(CLK), .RN(n695), .QN(n619) );
  DFFR_X1 REGISTERS_reg_20__24_ ( .D(n2946), .CK(CLK), .RN(n695), .QN(n620) );
  DFFR_X1 REGISTERS_reg_9__31_ ( .D(n3305), .CK(CLK), .RN(n610), .QN(n261) );
  DFFR_X1 REGISTERS_reg_9__30_ ( .D(n3304), .CK(CLK), .RN(n610), .QN(n262) );
  DFFR_X1 REGISTERS_reg_9__29_ ( .D(n3303), .CK(CLK), .RN(n610), .QN(n263) );
  DFFR_X1 REGISTERS_reg_9__28_ ( .D(n3302), .CK(CLK), .RN(n610), .QN(n264) );
  DFFR_X1 REGISTERS_reg_9__27_ ( .D(n3301), .CK(CLK), .RN(n610), .QN(n265) );
  DFFR_X1 REGISTERS_reg_9__26_ ( .D(n3300), .CK(CLK), .RN(n610), .QN(n266) );
  DFFR_X1 REGISTERS_reg_9__25_ ( .D(n3299), .CK(CLK), .RN(n610), .QN(n267) );
  DFFR_X1 REGISTERS_reg_9__24_ ( .D(n3298), .CK(CLK), .RN(n610), .QN(n268) );
  DFFR_X1 REGISTERS_reg_17__31_ ( .D(n3049), .CK(CLK), .RN(n704), .QN(n517) );
  DFFR_X1 REGISTERS_reg_17__30_ ( .D(n3048), .CK(CLK), .RN(n704), .QN(n518) );
  DFFR_X1 REGISTERS_reg_17__29_ ( .D(n3047), .CK(CLK), .RN(n703), .QN(n519) );
  DFFR_X1 REGISTERS_reg_17__28_ ( .D(n3046), .CK(CLK), .RN(n703), .QN(n520) );
  DFFR_X1 REGISTERS_reg_17__27_ ( .D(n3045), .CK(CLK), .RN(n703), .QN(n521) );
  DFFR_X1 REGISTERS_reg_17__26_ ( .D(n3044), .CK(CLK), .RN(n703), .QN(n522) );
  DFFR_X1 REGISTERS_reg_17__25_ ( .D(n3043), .CK(CLK), .RN(n703), .QN(n523) );
  DFFR_X1 REGISTERS_reg_17__24_ ( .D(n3042), .CK(CLK), .RN(n703), .QN(n524) );
  DFFR_X1 REGISTERS_reg_8__31_ ( .D(n3337), .CK(CLK), .RN(n666), .QN(n229) );
  DFFR_X1 REGISTERS_reg_8__30_ ( .D(n3336), .CK(CLK), .RN(n665), .QN(n230) );
  DFFR_X1 REGISTERS_reg_8__29_ ( .D(n3335), .CK(CLK), .RN(n665), .QN(n231) );
  DFFR_X1 REGISTERS_reg_8__28_ ( .D(n3334), .CK(CLK), .RN(n665), .QN(n232) );
  DFFR_X1 REGISTERS_reg_8__27_ ( .D(n3333), .CK(CLK), .RN(n665), .QN(n233) );
  DFFR_X1 REGISTERS_reg_8__26_ ( .D(n3332), .CK(CLK), .RN(n665), .QN(n234) );
  DFFR_X1 REGISTERS_reg_8__25_ ( .D(n3331), .CK(CLK), .RN(n665), .QN(n235) );
  DFFR_X1 REGISTERS_reg_8__24_ ( .D(n3330), .CK(CLK), .RN(n665), .QN(n236) );
  DFFR_X1 REGISTERS_reg_30__31_ ( .D(n2633), .CK(CLK), .RN(n690), .QN(n933) );
  DFFR_X1 REGISTERS_reg_30__30_ ( .D(n2632), .CK(CLK), .RN(n689), .QN(n934) );
  DFFR_X1 REGISTERS_reg_30__29_ ( .D(n2631), .CK(CLK), .RN(n689), .QN(n935) );
  DFFR_X1 REGISTERS_reg_30__28_ ( .D(n2630), .CK(CLK), .RN(n689), .QN(n936) );
  DFFR_X1 REGISTERS_reg_30__27_ ( .D(n2629), .CK(CLK), .RN(n689), .QN(n937) );
  DFFR_X1 REGISTERS_reg_30__26_ ( .D(n2628), .CK(CLK), .RN(n689), .QN(n938) );
  DFFR_X1 REGISTERS_reg_30__25_ ( .D(n2627), .CK(CLK), .RN(n689), .QN(n939) );
  DFFR_X1 REGISTERS_reg_30__24_ ( .D(n2626), .CK(CLK), .RN(n689), .QN(n940) );
  DFFR_X1 REGISTERS_reg_27__31_ ( .D(n2729), .CK(CLK), .RN(n677), .QN(n837) );
  DFFR_X1 REGISTERS_reg_27__30_ ( .D(n2728), .CK(CLK), .RN(n677), .QN(n838) );
  DFFR_X1 REGISTERS_reg_27__29_ ( .D(n2727), .CK(CLK), .RN(n677), .QN(n839) );
  DFFR_X1 REGISTERS_reg_27__28_ ( .D(n2726), .CK(CLK), .RN(n677), .QN(n840) );
  DFFR_X1 REGISTERS_reg_27__27_ ( .D(n2725), .CK(CLK), .RN(n676), .QN(n841) );
  DFFR_X1 REGISTERS_reg_27__26_ ( .D(n2724), .CK(CLK), .RN(n676), .QN(n842) );
  DFFR_X1 REGISTERS_reg_27__25_ ( .D(n2723), .CK(CLK), .RN(n676), .QN(n843) );
  DFFR_X1 REGISTERS_reg_27__24_ ( .D(n2722), .CK(CLK), .RN(n676), .QN(n844) );
  DFFR_X1 REGISTERS_reg_21__23_ ( .D(n2913), .CK(CLK), .RN(n713), .Q(n1157) );
  DFFR_X1 REGISTERS_reg_21__22_ ( .D(n2912), .CK(CLK), .RN(n713), .Q(n1158) );
  DFFR_X1 REGISTERS_reg_21__21_ ( .D(n2911), .CK(CLK), .RN(n713), .Q(n1159) );
  DFFR_X1 REGISTERS_reg_21__20_ ( .D(n2910), .CK(CLK), .RN(n713), .Q(n1160) );
  DFFR_X1 REGISTERS_reg_21__19_ ( .D(n2909), .CK(CLK), .RN(n713), .Q(n1161) );
  DFFR_X1 REGISTERS_reg_21__18_ ( .D(n2908), .CK(CLK), .RN(n712), .Q(n1162) );
  DFFR_X1 REGISTERS_reg_21__17_ ( .D(n2907), .CK(CLK), .RN(n712), .Q(n1163) );
  DFFR_X1 REGISTERS_reg_21__16_ ( .D(n2906), .CK(CLK), .RN(n712), .Q(n1164) );
  DFFR_X1 REGISTERS_reg_21__15_ ( .D(n2905), .CK(CLK), .RN(n712), .Q(n1165) );
  DFFR_X1 REGISTERS_reg_21__14_ ( .D(n2904), .CK(CLK), .RN(n712), .Q(n1166) );
  DFFR_X1 REGISTERS_reg_21__13_ ( .D(n2903), .CK(CLK), .RN(n712), .Q(n1167) );
  DFFR_X1 REGISTERS_reg_21__12_ ( .D(n2902), .CK(CLK), .RN(n712), .Q(n1168) );
  DFFR_X1 REGISTERS_reg_21__11_ ( .D(n2901), .CK(CLK), .RN(n712), .Q(n1169) );
  DFFR_X1 REGISTERS_reg_21__10_ ( .D(n2900), .CK(CLK), .RN(n712), .Q(n1170) );
  DFFR_X1 REGISTERS_reg_21__9_ ( .D(n2899), .CK(CLK), .RN(n712), .Q(n1171) );
  DFFR_X1 REGISTERS_reg_21__8_ ( .D(n2898), .CK(CLK), .RN(n712), .Q(n1172) );
  DFFR_X1 REGISTERS_reg_21__7_ ( .D(n2897), .CK(CLK), .RN(n712), .Q(n1173) );
  DFFR_X1 REGISTERS_reg_21__6_ ( .D(n2896), .CK(CLK), .RN(n711), .Q(n1174) );
  DFFR_X1 REGISTERS_reg_21__5_ ( .D(n2895), .CK(CLK), .RN(n711), .Q(n1175) );
  DFFR_X1 REGISTERS_reg_21__4_ ( .D(n2894), .CK(CLK), .RN(n711), .Q(n1176) );
  DFFR_X1 REGISTERS_reg_21__3_ ( .D(n2893), .CK(CLK), .RN(n711), .Q(n1177) );
  DFFR_X1 REGISTERS_reg_21__2_ ( .D(n2892), .CK(CLK), .RN(n711), .Q(n1178) );
  DFFR_X1 REGISTERS_reg_21__1_ ( .D(n2891), .CK(CLK), .RN(n711), .Q(n1179) );
  DFFR_X1 REGISTERS_reg_21__0_ ( .D(n2890), .CK(CLK), .RN(n711), .Q(n1180) );
  DFFR_X1 REGISTERS_reg_16__23_ ( .D(n3073), .CK(CLK), .RN(n611), .Q(n1055) );
  DFFR_X1 REGISTERS_reg_16__22_ ( .D(n3072), .CK(CLK), .RN(n611), .Q(n1056) );
  DFFR_X1 REGISTERS_reg_16__21_ ( .D(n3071), .CK(CLK), .RN(n611), .Q(n1057) );
  DFFR_X1 REGISTERS_reg_16__20_ ( .D(n3070), .CK(CLK), .RN(n611), .Q(n1058) );
  DFFR_X1 REGISTERS_reg_16__19_ ( .D(n3069), .CK(CLK), .RN(n611), .Q(n1059) );
  DFFR_X1 REGISTERS_reg_16__18_ ( .D(n3068), .CK(CLK), .RN(n611), .Q(n1060) );
  DFFR_X1 REGISTERS_reg_16__17_ ( .D(n3067), .CK(CLK), .RN(n611), .Q(n1061) );
  DFFR_X1 REGISTERS_reg_16__16_ ( .D(n3066), .CK(CLK), .RN(n648), .Q(n1062) );
  DFFR_X1 REGISTERS_reg_16__15_ ( .D(n3065), .CK(CLK), .RN(n653), .Q(n1063) );
  DFFR_X1 REGISTERS_reg_16__14_ ( .D(n3064), .CK(CLK), .RN(n705), .Q(n1064) );
  DFFR_X1 REGISTERS_reg_16__13_ ( .D(n3063), .CK(CLK), .RN(n705), .Q(n1065) );
  DFFR_X1 REGISTERS_reg_16__12_ ( .D(n3062), .CK(CLK), .RN(n705), .Q(n1066) );
  DFFR_X1 REGISTERS_reg_16__11_ ( .D(n3061), .CK(CLK), .RN(n705), .Q(n1067) );
  DFFR_X1 REGISTERS_reg_16__10_ ( .D(n3060), .CK(CLK), .RN(n705), .Q(n1068) );
  DFFR_X1 REGISTERS_reg_16__9_ ( .D(n3059), .CK(CLK), .RN(n704), .Q(n1069) );
  DFFR_X1 REGISTERS_reg_16__8_ ( .D(n3058), .CK(CLK), .RN(n704), .Q(n1070) );
  DFFR_X1 REGISTERS_reg_16__7_ ( .D(n3057), .CK(CLK), .RN(n704), .Q(n1071) );
  DFFR_X1 REGISTERS_reg_16__6_ ( .D(n3056), .CK(CLK), .RN(n704), .Q(n1072) );
  DFFR_X1 REGISTERS_reg_16__5_ ( .D(n3055), .CK(CLK), .RN(n704), .Q(n1073) );
  DFFR_X1 REGISTERS_reg_16__4_ ( .D(n3054), .CK(CLK), .RN(n704), .Q(n1074) );
  DFFR_X1 REGISTERS_reg_16__3_ ( .D(n3053), .CK(CLK), .RN(n704), .Q(n1075) );
  DFFR_X1 REGISTERS_reg_16__2_ ( .D(n3052), .CK(CLK), .RN(n704), .Q(n1076) );
  DFFR_X1 REGISTERS_reg_16__1_ ( .D(n3051), .CK(CLK), .RN(n704), .Q(n1077) );
  DFFR_X1 REGISTERS_reg_16__0_ ( .D(n3050), .CK(CLK), .RN(n704), .Q(n1078) );
  DFFR_X1 REGISTERS_reg_31__23_ ( .D(n2593), .CK(CLK), .RN(n686), .Q(n1298) );
  DFFR_X1 REGISTERS_reg_31__22_ ( .D(n2592), .CK(CLK), .RN(n686), .Q(n1299) );
  DFFR_X1 REGISTERS_reg_31__21_ ( .D(n2591), .CK(CLK), .RN(n686), .Q(n1300) );
  DFFR_X1 REGISTERS_reg_31__20_ ( .D(n2590), .CK(CLK), .RN(n686), .Q(n1301) );
  DFFR_X1 REGISTERS_reg_31__19_ ( .D(n2589), .CK(CLK), .RN(n686), .Q(n1302) );
  DFFR_X1 REGISTERS_reg_31__18_ ( .D(n2588), .CK(CLK), .RN(n686), .Q(n1303) );
  DFFR_X1 REGISTERS_reg_31__17_ ( .D(n2587), .CK(CLK), .RN(n686), .Q(n1304) );
  DFFR_X1 REGISTERS_reg_31__16_ ( .D(n2586), .CK(CLK), .RN(n686), .Q(n1305) );
  DFFR_X1 REGISTERS_reg_31__15_ ( .D(n2585), .CK(CLK), .RN(n685), .Q(n1306) );
  DFFR_X1 REGISTERS_reg_31__14_ ( .D(n2584), .CK(CLK), .RN(n685), .Q(n1307) );
  DFFR_X1 REGISTERS_reg_31__13_ ( .D(n2583), .CK(CLK), .RN(n685), .Q(n1308) );
  DFFR_X1 REGISTERS_reg_31__12_ ( .D(n2582), .CK(CLK), .RN(n685), .Q(n1309) );
  DFFR_X1 REGISTERS_reg_31__11_ ( .D(n2581), .CK(CLK), .RN(n685), .Q(n1310) );
  DFFR_X1 REGISTERS_reg_31__10_ ( .D(n2580), .CK(CLK), .RN(n685), .Q(n1311) );
  DFFR_X1 REGISTERS_reg_31__9_ ( .D(n2579), .CK(CLK), .RN(n685), .Q(n1312) );
  DFFR_X1 REGISTERS_reg_31__8_ ( .D(n2578), .CK(CLK), .RN(n685), .Q(n1313) );
  DFFR_X1 REGISTERS_reg_31__7_ ( .D(n2577), .CK(CLK), .RN(n685), .Q(n1314) );
  DFFR_X1 REGISTERS_reg_31__6_ ( .D(n2576), .CK(CLK), .RN(n685), .Q(n1315) );
  DFFR_X1 REGISTERS_reg_31__5_ ( .D(n2575), .CK(CLK), .RN(n685), .Q(n1316) );
  DFFR_X1 REGISTERS_reg_31__4_ ( .D(n2574), .CK(CLK), .RN(n685), .Q(n1317) );
  DFFR_X1 REGISTERS_reg_31__3_ ( .D(n2573), .CK(CLK), .RN(n684), .Q(n1318) );
  DFFR_X1 REGISTERS_reg_31__2_ ( .D(n2572), .CK(CLK), .RN(n684), .Q(n1319) );
  DFFR_X1 REGISTERS_reg_31__1_ ( .D(n2571), .CK(CLK), .RN(n684), .Q(n1320) );
  DFFR_X1 REGISTERS_reg_31__0_ ( .D(n2570), .CK(CLK), .RN(n689), .Q(n1321) );
  DFFR_X1 REGISTERS_reg_26__23_ ( .D(n2753), .CK(CLK), .RN(n679), .Q(n1196) );
  DFFR_X1 REGISTERS_reg_26__22_ ( .D(n2752), .CK(CLK), .RN(n679), .Q(n1197) );
  DFFR_X1 REGISTERS_reg_26__21_ ( .D(n2751), .CK(CLK), .RN(n679), .Q(n1198) );
  DFFR_X1 REGISTERS_reg_26__20_ ( .D(n2750), .CK(CLK), .RN(n679), .Q(n1199) );
  DFFR_X1 REGISTERS_reg_26__19_ ( .D(n2749), .CK(CLK), .RN(n678), .Q(n1200) );
  DFFR_X1 REGISTERS_reg_26__18_ ( .D(n2748), .CK(CLK), .RN(n678), .Q(n1201) );
  DFFR_X1 REGISTERS_reg_26__17_ ( .D(n2747), .CK(CLK), .RN(n678), .Q(n1202) );
  DFFR_X1 REGISTERS_reg_26__16_ ( .D(n2746), .CK(CLK), .RN(n678), .Q(n1203) );
  DFFR_X1 REGISTERS_reg_26__15_ ( .D(n2745), .CK(CLK), .RN(n678), .Q(n1204) );
  DFFR_X1 REGISTERS_reg_26__14_ ( .D(n2744), .CK(CLK), .RN(n678), .Q(n1205) );
  DFFR_X1 REGISTERS_reg_26__13_ ( .D(n2743), .CK(CLK), .RN(n678), .Q(n1206) );
  DFFR_X1 REGISTERS_reg_26__12_ ( .D(n2742), .CK(CLK), .RN(n678), .Q(n1207) );
  DFFR_X1 REGISTERS_reg_26__11_ ( .D(n2741), .CK(CLK), .RN(n678), .Q(n1208) );
  DFFR_X1 REGISTERS_reg_26__10_ ( .D(n2740), .CK(CLK), .RN(n678), .Q(n1209) );
  DFFR_X1 REGISTERS_reg_26__9_ ( .D(n2739), .CK(CLK), .RN(n678), .Q(n1210) );
  DFFR_X1 REGISTERS_reg_26__8_ ( .D(n2738), .CK(CLK), .RN(n678), .Q(n1211) );
  DFFR_X1 REGISTERS_reg_26__7_ ( .D(n2737), .CK(CLK), .RN(n677), .Q(n1212) );
  DFFR_X1 REGISTERS_reg_26__6_ ( .D(n2736), .CK(CLK), .RN(n677), .Q(n1213) );
  DFFR_X1 REGISTERS_reg_26__5_ ( .D(n2735), .CK(CLK), .RN(n677), .Q(n1214) );
  DFFR_X1 REGISTERS_reg_26__4_ ( .D(n2734), .CK(CLK), .RN(n677), .Q(n1215) );
  DFFR_X1 REGISTERS_reg_26__3_ ( .D(n2733), .CK(CLK), .RN(n677), .Q(n1216) );
  DFFR_X1 REGISTERS_reg_26__2_ ( .D(n2732), .CK(CLK), .RN(n677), .Q(n1217) );
  DFFR_X1 REGISTERS_reg_26__1_ ( .D(n2731), .CK(CLK), .RN(n677), .Q(n1218) );
  DFFR_X1 REGISTERS_reg_26__0_ ( .D(n2730), .CK(CLK), .RN(n677), .Q(n1219) );
  DFFR_X1 REGISTERS_reg_13__23_ ( .D(n3169), .CK(CLK), .RN(n652), .QN(n397) );
  DFFR_X1 REGISTERS_reg_13__22_ ( .D(n3168), .CK(CLK), .RN(n651), .QN(n398) );
  DFFR_X1 REGISTERS_reg_13__21_ ( .D(n3167), .CK(CLK), .RN(n651), .QN(n399) );
  DFFR_X1 REGISTERS_reg_13__20_ ( .D(n3166), .CK(CLK), .RN(n651), .QN(n400) );
  DFFR_X1 REGISTERS_reg_13__19_ ( .D(n3165), .CK(CLK), .RN(n651), .QN(n401) );
  DFFR_X1 REGISTERS_reg_13__18_ ( .D(n3164), .CK(CLK), .RN(n651), .QN(n402) );
  DFFR_X1 REGISTERS_reg_13__17_ ( .D(n3163), .CK(CLK), .RN(n651), .QN(n403) );
  DFFR_X1 REGISTERS_reg_13__16_ ( .D(n3162), .CK(CLK), .RN(n651), .QN(n404) );
  DFFR_X1 REGISTERS_reg_13__15_ ( .D(n3161), .CK(CLK), .RN(n651), .QN(n405) );
  DFFR_X1 REGISTERS_reg_13__14_ ( .D(n3160), .CK(CLK), .RN(n651), .QN(n406) );
  DFFR_X1 REGISTERS_reg_13__13_ ( .D(n3159), .CK(CLK), .RN(n651), .QN(n407) );
  DFFR_X1 REGISTERS_reg_13__12_ ( .D(n3158), .CK(CLK), .RN(n651), .QN(n408) );
  DFFR_X1 REGISTERS_reg_13__11_ ( .D(n3157), .CK(CLK), .RN(n651), .QN(n409) );
  DFFR_X1 REGISTERS_reg_13__10_ ( .D(n3156), .CK(CLK), .RN(n650), .QN(n410) );
  DFFR_X1 REGISTERS_reg_13__9_ ( .D(n3155), .CK(CLK), .RN(n650), .QN(n411) );
  DFFR_X1 REGISTERS_reg_13__8_ ( .D(n3154), .CK(CLK), .RN(n650), .QN(n412) );
  DFFR_X1 REGISTERS_reg_13__7_ ( .D(n3153), .CK(CLK), .RN(n650), .QN(n413) );
  DFFR_X1 REGISTERS_reg_13__6_ ( .D(n3152), .CK(CLK), .RN(n650), .QN(n414) );
  DFFR_X1 REGISTERS_reg_13__5_ ( .D(n3151), .CK(CLK), .RN(n650), .QN(n415) );
  DFFR_X1 REGISTERS_reg_13__4_ ( .D(n3150), .CK(CLK), .RN(n650), .QN(n416) );
  DFFR_X1 REGISTERS_reg_13__3_ ( .D(n3149), .CK(CLK), .RN(n650), .QN(n417) );
  DFFR_X1 REGISTERS_reg_13__2_ ( .D(n3148), .CK(CLK), .RN(n650), .QN(n418) );
  DFFR_X1 REGISTERS_reg_13__1_ ( .D(n3147), .CK(CLK), .RN(n650), .QN(n419) );
  DFFR_X1 REGISTERS_reg_13__0_ ( .D(n3146), .CK(CLK), .RN(n650), .QN(n420) );
  DFFR_X1 REGISTERS_reg_12__23_ ( .D(n3201), .CK(CLK), .RN(n602), .QN(n365) );
  DFFR_X1 REGISTERS_reg_12__22_ ( .D(n3200), .CK(CLK), .RN(n601), .QN(n366) );
  DFFR_X1 REGISTERS_reg_12__21_ ( .D(n3199), .CK(CLK), .RN(n601), .QN(n367) );
  DFFR_X1 REGISTERS_reg_12__20_ ( .D(n3198), .CK(CLK), .RN(n601), .QN(n368) );
  DFFR_X1 REGISTERS_reg_12__19_ ( .D(n3197), .CK(CLK), .RN(n601), .QN(n369) );
  DFFR_X1 REGISTERS_reg_12__18_ ( .D(n3196), .CK(CLK), .RN(n601), .QN(n370) );
  DFFR_X1 REGISTERS_reg_12__17_ ( .D(n3195), .CK(CLK), .RN(n601), .QN(n371) );
  DFFR_X1 REGISTERS_reg_12__16_ ( .D(n3194), .CK(CLK), .RN(n601), .QN(n372) );
  DFFR_X1 REGISTERS_reg_12__15_ ( .D(n3193), .CK(CLK), .RN(n601), .QN(n373) );
  DFFR_X1 REGISTERS_reg_7__31_ ( .D(n3369), .CK(CLK), .RN(n668), .Q(n4350), 
        .QN(n1374) );
  DFFR_X1 REGISTERS_reg_7__30_ ( .D(n3368), .CK(CLK), .RN(n668), .Q(n4349), 
        .QN(n1404) );
  DFFR_X1 REGISTERS_reg_7__29_ ( .D(n3367), .CK(CLK), .RN(n668), .Q(n4348), 
        .QN(n1429) );
  DFFR_X1 REGISTERS_reg_7__28_ ( .D(n3366), .CK(CLK), .RN(n668), .Q(n4347), 
        .QN(n1454) );
  DFFR_X1 REGISTERS_reg_7__27_ ( .D(n3365), .CK(CLK), .RN(n668), .Q(n4346), 
        .QN(n1479) );
  DFFR_X1 REGISTERS_reg_7__26_ ( .D(n3364), .CK(CLK), .RN(n668), .Q(n4345), 
        .QN(n1504) );
  DFFR_X1 REGISTERS_reg_7__25_ ( .D(n3363), .CK(CLK), .RN(n668), .Q(n4344), 
        .QN(n1529) );
  DFFR_X1 REGISTERS_reg_7__24_ ( .D(n3362), .CK(CLK), .RN(n668), .Q(n4343), 
        .QN(n1554) );
  DFFR_X1 REGISTERS_reg_6__31_ ( .D(n3401), .CK(CLK), .RN(n671), .Q(n4382), 
        .QN(n1372) );
  DFFR_X1 REGISTERS_reg_6__30_ ( .D(n3400), .CK(CLK), .RN(n671), .Q(n4381), 
        .QN(n1403) );
  DFFR_X1 REGISTERS_reg_6__29_ ( .D(n3399), .CK(CLK), .RN(n671), .Q(n4380), 
        .QN(n1428) );
  DFFR_X1 REGISTERS_reg_6__28_ ( .D(n3398), .CK(CLK), .RN(n671), .Q(n4379), 
        .QN(n1453) );
  DFFR_X1 REGISTERS_reg_6__27_ ( .D(n3397), .CK(CLK), .RN(n671), .Q(n4378), 
        .QN(n1478) );
  DFFR_X1 REGISTERS_reg_6__26_ ( .D(n3396), .CK(CLK), .RN(n671), .Q(n4377), 
        .QN(n1503) );
  DFFR_X1 REGISTERS_reg_6__25_ ( .D(n3395), .CK(CLK), .RN(n670), .Q(n4376), 
        .QN(n1528) );
  DFFR_X1 REGISTERS_reg_6__24_ ( .D(n3394), .CK(CLK), .RN(n670), .Q(n4375), 
        .QN(n1553) );
  DFFR_X1 REGISTERS_reg_3__31_ ( .D(n3497), .CK(CLK), .RN(n658), .Q(n4414), 
        .QN(n1381) );
  DFFR_X1 REGISTERS_reg_3__30_ ( .D(n3496), .CK(CLK), .RN(n658), .Q(n4413), 
        .QN(n1407) );
  DFFR_X1 REGISTERS_reg_3__29_ ( .D(n3495), .CK(CLK), .RN(n658), .Q(n4412), 
        .QN(n1432) );
  DFFR_X1 REGISTERS_reg_3__28_ ( .D(n3494), .CK(CLK), .RN(n658), .Q(n4411), 
        .QN(n1457) );
  DFFR_X1 REGISTERS_reg_3__27_ ( .D(n3493), .CK(CLK), .RN(n658), .Q(n4410), 
        .QN(n1482) );
  DFFR_X1 REGISTERS_reg_3__26_ ( .D(n3492), .CK(CLK), .RN(n658), .Q(n4409), 
        .QN(n1507) );
  DFFR_X1 REGISTERS_reg_3__25_ ( .D(n3491), .CK(CLK), .RN(n658), .Q(n4408), 
        .QN(n1532) );
  DFFR_X1 REGISTERS_reg_3__24_ ( .D(n3490), .CK(CLK), .RN(n658), .Q(n4407), 
        .QN(n1557) );
  DFFR_X1 REGISTERS_reg_2__31_ ( .D(n3529), .CK(CLK), .RN(n661), .Q(n4446), 
        .QN(n1379) );
  DFFR_X1 REGISTERS_reg_2__30_ ( .D(n3528), .CK(CLK), .RN(n661), .Q(n4445), 
        .QN(n1406) );
  DFFR_X1 REGISTERS_reg_2__29_ ( .D(n3527), .CK(CLK), .RN(n661), .Q(n4444), 
        .QN(n1431) );
  DFFR_X1 REGISTERS_reg_2__28_ ( .D(n3526), .CK(CLK), .RN(n661), .Q(n4443), 
        .QN(n1456) );
  DFFR_X1 REGISTERS_reg_2__27_ ( .D(n3525), .CK(CLK), .RN(n661), .Q(n4442), 
        .QN(n1481) );
  DFFR_X1 REGISTERS_reg_2__26_ ( .D(n3524), .CK(CLK), .RN(n661), .Q(n4441), 
        .QN(n1506) );
  DFFR_X1 REGISTERS_reg_2__25_ ( .D(n3523), .CK(CLK), .RN(n661), .Q(n4440), 
        .QN(n1531) );
  DFFR_X1 REGISTERS_reg_2__24_ ( .D(n3522), .CK(CLK), .RN(n660), .Q(n4439), 
        .QN(n1556) );
  DFFR_X1 REGISTERS_reg_15__31_ ( .D(n3113), .CK(CLK), .RN(n647), .Q(n4222) );
  DFFR_X1 REGISTERS_reg_15__30_ ( .D(n3112), .CK(CLK), .RN(n647), .Q(n4221) );
  DFFR_X1 REGISTERS_reg_15__29_ ( .D(n3111), .CK(CLK), .RN(n647), .Q(n4220) );
  DFFR_X1 REGISTERS_reg_15__28_ ( .D(n3110), .CK(CLK), .RN(n647), .Q(n4219) );
  DFFR_X1 REGISTERS_reg_15__27_ ( .D(n3109), .CK(CLK), .RN(n646), .Q(n4218) );
  DFFR_X1 REGISTERS_reg_15__26_ ( .D(n3108), .CK(CLK), .RN(n646), .Q(n4217) );
  DFFR_X1 REGISTERS_reg_15__25_ ( .D(n3107), .CK(CLK), .RN(n646), .Q(n4216) );
  DFFR_X1 REGISTERS_reg_15__24_ ( .D(n3106), .CK(CLK), .RN(n646), .Q(n4215) );
  DFFR_X1 REGISTERS_reg_14__31_ ( .D(n3145), .CK(CLK), .RN(n650), .Q(n4254) );
  DFFR_X1 REGISTERS_reg_14__30_ ( .D(n3144), .CK(CLK), .RN(n649), .Q(n4253) );
  DFFR_X1 REGISTERS_reg_14__29_ ( .D(n3143), .CK(CLK), .RN(n649), .Q(n4252) );
  DFFR_X1 REGISTERS_reg_14__28_ ( .D(n3142), .CK(CLK), .RN(n649), .Q(n4251) );
  DFFR_X1 REGISTERS_reg_14__27_ ( .D(n3141), .CK(CLK), .RN(n649), .Q(n4250) );
  DFFR_X1 REGISTERS_reg_14__26_ ( .D(n3140), .CK(CLK), .RN(n649), .Q(n4249) );
  DFFR_X1 REGISTERS_reg_14__25_ ( .D(n3139), .CK(CLK), .RN(n649), .Q(n4248) );
  DFFR_X1 REGISTERS_reg_14__24_ ( .D(n3138), .CK(CLK), .RN(n649), .Q(n4247) );
  DFFR_X1 REGISTERS_reg_23__31_ ( .D(n2857), .CK(CLK), .RN(n708), .Q(n4094), 
        .QN(n1333) );
  DFFR_X1 REGISTERS_reg_23__30_ ( .D(n2856), .CK(CLK), .RN(n708), .Q(n4093), 
        .QN(n1388) );
  DFFR_X1 REGISTERS_reg_23__29_ ( .D(n2855), .CK(CLK), .RN(n708), .Q(n4092), 
        .QN(n1413) );
  DFFR_X1 REGISTERS_reg_23__28_ ( .D(n2854), .CK(CLK), .RN(n708), .Q(n4091), 
        .QN(n1438) );
  DFFR_X1 REGISTERS_reg_23__27_ ( .D(n2853), .CK(CLK), .RN(n708), .Q(n4090), 
        .QN(n1463) );
  DFFR_X1 REGISTERS_reg_23__26_ ( .D(n2852), .CK(CLK), .RN(n708), .Q(n4089), 
        .QN(n1488) );
  DFFR_X1 REGISTERS_reg_23__25_ ( .D(n2851), .CK(CLK), .RN(n708), .Q(n4088), 
        .QN(n1513) );
  DFFR_X1 REGISTERS_reg_23__24_ ( .D(n2850), .CK(CLK), .RN(n708), .Q(n4087), 
        .QN(n1538) );
  DFFR_X1 REGISTERS_reg_22__31_ ( .D(n2889), .CK(CLK), .RN(n711), .Q(n4126), 
        .QN(n1351) );
  DFFR_X1 REGISTERS_reg_22__30_ ( .D(n2888), .CK(CLK), .RN(n711), .Q(n4125), 
        .QN(n1395) );
  DFFR_X1 REGISTERS_reg_22__29_ ( .D(n2887), .CK(CLK), .RN(n711), .Q(n4124), 
        .QN(n1420) );
  DFFR_X1 REGISTERS_reg_22__28_ ( .D(n2886), .CK(CLK), .RN(n711), .Q(n4123), 
        .QN(n1445) );
  DFFR_X1 REGISTERS_reg_22__27_ ( .D(n2885), .CK(CLK), .RN(n711), .Q(n4122), 
        .QN(n1470) );
  DFFR_X1 REGISTERS_reg_22__26_ ( .D(n2884), .CK(CLK), .RN(n710), .Q(n4121), 
        .QN(n1495) );
  DFFR_X1 REGISTERS_reg_22__25_ ( .D(n2883), .CK(CLK), .RN(n710), .Q(n4120), 
        .QN(n1520) );
  DFFR_X1 REGISTERS_reg_22__24_ ( .D(n2882), .CK(CLK), .RN(n710), .Q(n4119), 
        .QN(n1545) );
  DFFR_X1 REGISTERS_reg_11__31_ ( .D(n3241), .CK(CLK), .RN(n605), .Q(n4286) );
  DFFR_X1 REGISTERS_reg_11__30_ ( .D(n3240), .CK(CLK), .RN(n605), .Q(n4285) );
  DFFR_X1 REGISTERS_reg_11__29_ ( .D(n3239), .CK(CLK), .RN(n605), .Q(n4284) );
  DFFR_X1 REGISTERS_reg_11__28_ ( .D(n3238), .CK(CLK), .RN(n605), .Q(n4283) );
  DFFR_X1 REGISTERS_reg_11__27_ ( .D(n3237), .CK(CLK), .RN(n605), .Q(n4282) );
  DFFR_X1 REGISTERS_reg_11__26_ ( .D(n3236), .CK(CLK), .RN(n604), .Q(n4281) );
  DFFR_X1 REGISTERS_reg_11__25_ ( .D(n3235), .CK(CLK), .RN(n604), .Q(n4280) );
  DFFR_X1 REGISTERS_reg_11__24_ ( .D(n3234), .CK(CLK), .RN(n604), .Q(n4279) );
  DFFR_X1 REGISTERS_reg_10__31_ ( .D(n3273), .CK(CLK), .RN(n608), .Q(n4318) );
  DFFR_X1 REGISTERS_reg_10__30_ ( .D(n3272), .CK(CLK), .RN(n608), .Q(n4317) );
  DFFR_X1 REGISTERS_reg_10__29_ ( .D(n3271), .CK(CLK), .RN(n607), .Q(n4316) );
  DFFR_X1 REGISTERS_reg_10__28_ ( .D(n3270), .CK(CLK), .RN(n607), .Q(n4315) );
  DFFR_X1 REGISTERS_reg_10__27_ ( .D(n3269), .CK(CLK), .RN(n607), .Q(n4314) );
  DFFR_X1 REGISTERS_reg_10__26_ ( .D(n3268), .CK(CLK), .RN(n607), .Q(n4313) );
  DFFR_X1 REGISTERS_reg_10__25_ ( .D(n3267), .CK(CLK), .RN(n607), .Q(n4312) );
  DFFR_X1 REGISTERS_reg_10__24_ ( .D(n3266), .CK(CLK), .RN(n607), .Q(n4311) );
  DFFR_X1 REGISTERS_reg_19__31_ ( .D(n2985), .CK(CLK), .RN(n698), .Q(n4158) );
  DFFR_X1 REGISTERS_reg_19__30_ ( .D(n2984), .CK(CLK), .RN(n698), .Q(n4157) );
  DFFR_X1 REGISTERS_reg_19__29_ ( .D(n2983), .CK(CLK), .RN(n698), .Q(n4156) );
  DFFR_X1 REGISTERS_reg_19__28_ ( .D(n2982), .CK(CLK), .RN(n698), .Q(n4155) );
  DFFR_X1 REGISTERS_reg_19__27_ ( .D(n2981), .CK(CLK), .RN(n698), .Q(n4154) );
  DFFR_X1 REGISTERS_reg_19__26_ ( .D(n2980), .CK(CLK), .RN(n698), .Q(n4153) );
  DFFR_X1 REGISTERS_reg_19__25_ ( .D(n2979), .CK(CLK), .RN(n698), .Q(n4152) );
  DFFR_X1 REGISTERS_reg_19__24_ ( .D(n2978), .CK(CLK), .RN(n698), .Q(n4151) );
  DFFR_X1 REGISTERS_reg_18__31_ ( .D(n3017), .CK(CLK), .RN(n701), .Q(n4190) );
  DFFR_X1 REGISTERS_reg_18__30_ ( .D(n3016), .CK(CLK), .RN(n701), .Q(n4189) );
  DFFR_X1 REGISTERS_reg_18__29_ ( .D(n3015), .CK(CLK), .RN(n701), .Q(n4188) );
  DFFR_X1 REGISTERS_reg_18__28_ ( .D(n3014), .CK(CLK), .RN(n701), .Q(n4187) );
  DFFR_X1 REGISTERS_reg_18__27_ ( .D(n3013), .CK(CLK), .RN(n701), .Q(n4186) );
  DFFR_X1 REGISTERS_reg_18__26_ ( .D(n3012), .CK(CLK), .RN(n701), .Q(n4185) );
  DFFR_X1 REGISTERS_reg_18__25_ ( .D(n3011), .CK(CLK), .RN(n700), .Q(n4184) );
  DFFR_X1 REGISTERS_reg_18__24_ ( .D(n3010), .CK(CLK), .RN(n700), .Q(n4183) );
  DFFR_X1 REGISTERS_reg_29__31_ ( .D(n2665), .CK(CLK), .RN(n692), .Q(n3966) );
  DFFR_X1 REGISTERS_reg_29__30_ ( .D(n2664), .CK(CLK), .RN(n692), .Q(n3965) );
  DFFR_X1 REGISTERS_reg_29__29_ ( .D(n2663), .CK(CLK), .RN(n692), .Q(n3964) );
  DFFR_X1 REGISTERS_reg_29__28_ ( .D(n2662), .CK(CLK), .RN(n692), .Q(n3963) );
  DFFR_X1 REGISTERS_reg_29__27_ ( .D(n2661), .CK(CLK), .RN(n692), .Q(n3962) );
  DFFR_X1 REGISTERS_reg_29__26_ ( .D(n2660), .CK(CLK), .RN(n692), .Q(n3961) );
  DFFR_X1 REGISTERS_reg_29__25_ ( .D(n2659), .CK(CLK), .RN(n692), .Q(n3960) );
  DFFR_X1 REGISTERS_reg_29__24_ ( .D(n2658), .CK(CLK), .RN(n692), .Q(n3959) );
  DFFR_X1 REGISTERS_reg_28__31_ ( .D(n2697), .CK(CLK), .RN(n674), .Q(n3998), 
        .QN(n1338) );
  DFFR_X1 REGISTERS_reg_28__30_ ( .D(n2696), .CK(CLK), .RN(n674), .Q(n3997), 
        .QN(n1390) );
  DFFR_X1 REGISTERS_reg_28__29_ ( .D(n2695), .CK(CLK), .RN(n674), .Q(n3996), 
        .QN(n1415) );
  DFFR_X1 REGISTERS_reg_28__28_ ( .D(n2694), .CK(CLK), .RN(n679), .Q(n3995), 
        .QN(n1440) );
  DFFR_X1 REGISTERS_reg_28__27_ ( .D(n2693), .CK(CLK), .RN(n694), .Q(n3994), 
        .QN(n1465) );
  DFFR_X1 REGISTERS_reg_28__26_ ( .D(n2692), .CK(CLK), .RN(n695), .Q(n3993), 
        .QN(n1490) );
  DFFR_X1 REGISTERS_reg_28__25_ ( .D(n2691), .CK(CLK), .RN(n694), .Q(n3992), 
        .QN(n1515) );
  DFFR_X1 REGISTERS_reg_28__24_ ( .D(n2690), .CK(CLK), .RN(n694), .Q(n3991), 
        .QN(n1540) );
  DFFR_X1 REGISTERS_reg_25__31_ ( .D(n2793), .CK(CLK), .RN(n682), .Q(n4030) );
  DFFR_X1 REGISTERS_reg_25__30_ ( .D(n2792), .CK(CLK), .RN(n682), .Q(n4029) );
  DFFR_X1 REGISTERS_reg_25__29_ ( .D(n2791), .CK(CLK), .RN(n682), .Q(n4028) );
  DFFR_X1 REGISTERS_reg_25__28_ ( .D(n2790), .CK(CLK), .RN(n682), .Q(n4027) );
  DFFR_X1 REGISTERS_reg_25__27_ ( .D(n2789), .CK(CLK), .RN(n682), .Q(n4026) );
  DFFR_X1 REGISTERS_reg_25__26_ ( .D(n2788), .CK(CLK), .RN(n682), .Q(n4025) );
  DFFR_X1 REGISTERS_reg_25__25_ ( .D(n2787), .CK(CLK), .RN(n682), .Q(n4024) );
  DFFR_X1 REGISTERS_reg_25__24_ ( .D(n2786), .CK(CLK), .RN(n682), .Q(n4023) );
  DFFR_X1 REGISTERS_reg_24__31_ ( .D(n2825), .CK(CLK), .RN(n705), .Q(n4062) );
  DFFR_X1 REGISTERS_reg_24__30_ ( .D(n2824), .CK(CLK), .RN(n705), .Q(n4061) );
  DFFR_X1 REGISTERS_reg_24__29_ ( .D(n2823), .CK(CLK), .RN(n705), .Q(n4060) );
  DFFR_X1 REGISTERS_reg_24__28_ ( .D(n2822), .CK(CLK), .RN(n705), .Q(n4059) );
  DFFR_X1 REGISTERS_reg_24__27_ ( .D(n2821), .CK(CLK), .RN(n705), .Q(n4058) );
  DFFR_X1 REGISTERS_reg_24__26_ ( .D(n2820), .CK(CLK), .RN(n705), .Q(n4057) );
  DFFR_X1 REGISTERS_reg_24__25_ ( .D(n2819), .CK(CLK), .RN(n705), .Q(n4056) );
  DFFR_X1 REGISTERS_reg_24__24_ ( .D(n2818), .CK(CLK), .RN(n710), .Q(n4055) );
  DFFR_X1 REGISTERS_reg_7__23_ ( .D(n3361), .CK(CLK), .RN(n668), .Q(n4342), 
        .QN(n1579) );
  DFFR_X1 REGISTERS_reg_7__22_ ( .D(n3360), .CK(CLK), .RN(n667), .Q(n4341), 
        .QN(n1604) );
  DFFR_X1 REGISTERS_reg_7__21_ ( .D(n3359), .CK(CLK), .RN(n667), .Q(n4340), 
        .QN(n1629) );
  DFFR_X1 REGISTERS_reg_7__20_ ( .D(n3358), .CK(CLK), .RN(n667), .Q(n4339), 
        .QN(n1654) );
  DFFR_X1 REGISTERS_reg_7__19_ ( .D(n3357), .CK(CLK), .RN(n667), .Q(n4338), 
        .QN(n1679) );
  DFFR_X1 REGISTERS_reg_7__18_ ( .D(n3356), .CK(CLK), .RN(n667), .Q(n4337), 
        .QN(n1704) );
  DFFR_X1 REGISTERS_reg_7__17_ ( .D(n3355), .CK(CLK), .RN(n667), .Q(n4336), 
        .QN(n1729) );
  DFFR_X1 REGISTERS_reg_7__16_ ( .D(n3354), .CK(CLK), .RN(n667), .Q(n4335), 
        .QN(n1754) );
  DFFR_X1 REGISTERS_reg_7__15_ ( .D(n3353), .CK(CLK), .RN(n667), .Q(n4334), 
        .QN(n1779) );
  DFFR_X1 REGISTERS_reg_7__14_ ( .D(n3352), .CK(CLK), .RN(n667), .Q(n4333), 
        .QN(n1804) );
  DFFR_X1 REGISTERS_reg_7__13_ ( .D(n3351), .CK(CLK), .RN(n667), .Q(n4332), 
        .QN(n1829) );
  DFFR_X1 REGISTERS_reg_7__12_ ( .D(n3350), .CK(CLK), .RN(n667), .Q(n4331), 
        .QN(n1854) );
  DFFR_X1 REGISTERS_reg_7__11_ ( .D(n3349), .CK(CLK), .RN(n667), .Q(n4330), 
        .QN(n1879) );
  DFFR_X1 REGISTERS_reg_7__10_ ( .D(n3348), .CK(CLK), .RN(n666), .Q(n4329), 
        .QN(n1904) );
  DFFR_X1 REGISTERS_reg_7__9_ ( .D(n3347), .CK(CLK), .RN(n666), .Q(n4328), 
        .QN(n1929) );
  DFFR_X1 REGISTERS_reg_7__8_ ( .D(n3346), .CK(CLK), .RN(n666), .Q(n4327), 
        .QN(n1954) );
  DFFR_X1 REGISTERS_reg_7__7_ ( .D(n3345), .CK(CLK), .RN(n666), .Q(n4326), 
        .QN(n1979) );
  DFFR_X1 REGISTERS_reg_7__6_ ( .D(n3344), .CK(CLK), .RN(n666), .Q(n4325), 
        .QN(n2004) );
  DFFR_X1 REGISTERS_reg_7__5_ ( .D(n3343), .CK(CLK), .RN(n666), .Q(n4324), 
        .QN(n2029) );
  DFFR_X1 REGISTERS_reg_7__4_ ( .D(n3342), .CK(CLK), .RN(n666), .Q(n4323), 
        .QN(n2054) );
  DFFR_X1 REGISTERS_reg_7__3_ ( .D(n3341), .CK(CLK), .RN(n666), .Q(n4322), 
        .QN(n2079) );
  DFFR_X1 REGISTERS_reg_7__2_ ( .D(n3340), .CK(CLK), .RN(n666), .Q(n4321), 
        .QN(n2104) );
  DFFR_X1 REGISTERS_reg_7__1_ ( .D(n3339), .CK(CLK), .RN(n666), .Q(n4320), 
        .QN(n2129) );
  DFFR_X1 REGISTERS_reg_7__0_ ( .D(n3338), .CK(CLK), .RN(n666), .Q(n4319), 
        .QN(n2167) );
  DFFR_X1 REGISTERS_reg_6__23_ ( .D(n3393), .CK(CLK), .RN(n670), .Q(n4374), 
        .QN(n1578) );
  DFFR_X1 REGISTERS_reg_6__22_ ( .D(n3392), .CK(CLK), .RN(n670), .Q(n4373), 
        .QN(n1603) );
  DFFR_X1 REGISTERS_reg_6__21_ ( .D(n3391), .CK(CLK), .RN(n670), .Q(n4372), 
        .QN(n1628) );
  DFFR_X1 REGISTERS_reg_6__20_ ( .D(n3390), .CK(CLK), .RN(n670), .Q(n4371), 
        .QN(n1653) );
  DFFR_X1 REGISTERS_reg_6__19_ ( .D(n3389), .CK(CLK), .RN(n670), .Q(n4370), 
        .QN(n1678) );
  DFFR_X1 REGISTERS_reg_6__18_ ( .D(n3388), .CK(CLK), .RN(n670), .Q(n4369), 
        .QN(n1703) );
  DFFR_X1 REGISTERS_reg_6__17_ ( .D(n3387), .CK(CLK), .RN(n670), .Q(n4368), 
        .QN(n1728) );
  DFFR_X1 REGISTERS_reg_6__16_ ( .D(n3386), .CK(CLK), .RN(n670), .Q(n4367), 
        .QN(n1753) );
  DFFR_X1 REGISTERS_reg_6__15_ ( .D(n3385), .CK(CLK), .RN(n670), .Q(n4366), 
        .QN(n1778) );
  DFFR_X1 REGISTERS_reg_6__14_ ( .D(n3384), .CK(CLK), .RN(n670), .Q(n4365), 
        .QN(n1803) );
  DFFR_X1 REGISTERS_reg_6__13_ ( .D(n3383), .CK(CLK), .RN(n669), .Q(n4364), 
        .QN(n1828) );
  DFFR_X1 REGISTERS_reg_6__12_ ( .D(n3382), .CK(CLK), .RN(n669), .Q(n4363), 
        .QN(n1853) );
  DFFR_X1 REGISTERS_reg_6__11_ ( .D(n3381), .CK(CLK), .RN(n669), .Q(n4362), 
        .QN(n1878) );
  DFFR_X1 REGISTERS_reg_6__10_ ( .D(n3380), .CK(CLK), .RN(n669), .Q(n4361), 
        .QN(n1903) );
  DFFR_X1 REGISTERS_reg_6__9_ ( .D(n3379), .CK(CLK), .RN(n669), .Q(n4360), 
        .QN(n1928) );
  DFFR_X1 REGISTERS_reg_6__8_ ( .D(n3378), .CK(CLK), .RN(n669), .Q(n4359), 
        .QN(n1953) );
  DFFR_X1 REGISTERS_reg_6__7_ ( .D(n3377), .CK(CLK), .RN(n669), .Q(n4358), 
        .QN(n1978) );
  DFFR_X1 REGISTERS_reg_6__6_ ( .D(n3376), .CK(CLK), .RN(n669), .Q(n4357), 
        .QN(n2003) );
  DFFR_X1 REGISTERS_reg_6__5_ ( .D(n3375), .CK(CLK), .RN(n669), .Q(n4356), 
        .QN(n2028) );
  DFFR_X1 REGISTERS_reg_6__4_ ( .D(n3374), .CK(CLK), .RN(n669), .Q(n4355), 
        .QN(n2053) );
  DFFR_X1 REGISTERS_reg_6__3_ ( .D(n3373), .CK(CLK), .RN(n669), .Q(n4354), 
        .QN(n2078) );
  DFFR_X1 REGISTERS_reg_6__2_ ( .D(n3372), .CK(CLK), .RN(n668), .Q(n4353), 
        .QN(n2103) );
  DFFR_X1 REGISTERS_reg_6__1_ ( .D(n3371), .CK(CLK), .RN(n668), .Q(n4352), 
        .QN(n2128) );
  DFFR_X1 REGISTERS_reg_6__0_ ( .D(n3370), .CK(CLK), .RN(n668), .Q(n4351), 
        .QN(n2166) );
  DFFR_X1 REGISTERS_reg_3__23_ ( .D(n3489), .CK(CLK), .RN(n658), .Q(n4406), 
        .QN(n1582) );
  DFFR_X1 REGISTERS_reg_3__22_ ( .D(n3488), .CK(CLK), .RN(n658), .Q(n4405), 
        .QN(n1607) );
  DFFR_X1 REGISTERS_reg_3__21_ ( .D(n3487), .CK(CLK), .RN(n657), .Q(n4404), 
        .QN(n1632) );
  DFFR_X1 REGISTERS_reg_3__20_ ( .D(n3486), .CK(CLK), .RN(n657), .Q(n4403), 
        .QN(n1657) );
  DFFR_X1 REGISTERS_reg_3__19_ ( .D(n3485), .CK(CLK), .RN(n657), .Q(n4402), 
        .QN(n1682) );
  DFFR_X1 REGISTERS_reg_3__18_ ( .D(n3484), .CK(CLK), .RN(n657), .Q(n4401), 
        .QN(n1707) );
  DFFR_X1 REGISTERS_reg_3__17_ ( .D(n3483), .CK(CLK), .RN(n657), .Q(n4400), 
        .QN(n1732) );
  DFFR_X1 REGISTERS_reg_3__16_ ( .D(n3482), .CK(CLK), .RN(n657), .Q(n4399), 
        .QN(n1757) );
  DFFR_X1 REGISTERS_reg_3__15_ ( .D(n3481), .CK(CLK), .RN(n657), .Q(n4398), 
        .QN(n1782) );
  DFFR_X1 REGISTERS_reg_3__14_ ( .D(n3480), .CK(CLK), .RN(n657), .Q(n4397), 
        .QN(n1807) );
  DFFR_X1 REGISTERS_reg_3__13_ ( .D(n3479), .CK(CLK), .RN(n657), .Q(n4396), 
        .QN(n1832) );
  DFFR_X1 REGISTERS_reg_3__12_ ( .D(n3478), .CK(CLK), .RN(n657), .Q(n4395), 
        .QN(n1857) );
  DFFR_X1 REGISTERS_reg_3__11_ ( .D(n3477), .CK(CLK), .RN(n657), .Q(n4394), 
        .QN(n1882) );
  DFFR_X1 REGISTERS_reg_3__10_ ( .D(n3476), .CK(CLK), .RN(n657), .Q(n4393), 
        .QN(n1907) );
  DFFR_X1 REGISTERS_reg_3__9_ ( .D(n3475), .CK(CLK), .RN(n656), .Q(n4392), 
        .QN(n1932) );
  DFFR_X1 REGISTERS_reg_3__8_ ( .D(n3474), .CK(CLK), .RN(n656), .Q(n4391), 
        .QN(n1957) );
  DFFR_X1 REGISTERS_reg_3__7_ ( .D(n3473), .CK(CLK), .RN(n656), .Q(n4390), 
        .QN(n1982) );
  DFFR_X1 REGISTERS_reg_3__6_ ( .D(n3472), .CK(CLK), .RN(n656), .Q(n4389), 
        .QN(n2007) );
  DFFR_X1 REGISTERS_reg_3__5_ ( .D(n3471), .CK(CLK), .RN(n656), .Q(n4388), 
        .QN(n2032) );
  DFFR_X1 REGISTERS_reg_3__4_ ( .D(n3470), .CK(CLK), .RN(n656), .Q(n4387), 
        .QN(n2057) );
  DFFR_X1 REGISTERS_reg_3__3_ ( .D(n3469), .CK(CLK), .RN(n656), .Q(n4386), 
        .QN(n2082) );
  DFFR_X1 REGISTERS_reg_3__2_ ( .D(n3468), .CK(CLK), .RN(n656), .Q(n4385), 
        .QN(n2107) );
  DFFR_X1 REGISTERS_reg_3__1_ ( .D(n3467), .CK(CLK), .RN(n656), .Q(n4384), 
        .QN(n2132) );
  DFFR_X1 REGISTERS_reg_3__0_ ( .D(n3466), .CK(CLK), .RN(n656), .Q(n4383), 
        .QN(n2172) );
  DFFR_X1 REGISTERS_reg_2__23_ ( .D(n3521), .CK(CLK), .RN(n660), .Q(n4438), 
        .QN(n1581) );
  DFFR_X1 REGISTERS_reg_2__22_ ( .D(n3520), .CK(CLK), .RN(n660), .Q(n4437), 
        .QN(n1606) );
  DFFR_X1 REGISTERS_reg_2__21_ ( .D(n3519), .CK(CLK), .RN(n660), .Q(n4436), 
        .QN(n1631) );
  DFFR_X1 REGISTERS_reg_2__20_ ( .D(n3518), .CK(CLK), .RN(n660), .Q(n4435), 
        .QN(n1656) );
  DFFR_X1 REGISTERS_reg_2__19_ ( .D(n3517), .CK(CLK), .RN(n660), .Q(n4434), 
        .QN(n1681) );
  DFFR_X1 REGISTERS_reg_2__18_ ( .D(n3516), .CK(CLK), .RN(n660), .Q(n4433), 
        .QN(n1706) );
  DFFR_X1 REGISTERS_reg_2__17_ ( .D(n3515), .CK(CLK), .RN(n660), .Q(n4432), 
        .QN(n1731) );
  DFFR_X1 REGISTERS_reg_2__16_ ( .D(n3514), .CK(CLK), .RN(n660), .Q(n4431), 
        .QN(n1756) );
  DFFR_X1 REGISTERS_reg_2__15_ ( .D(n3513), .CK(CLK), .RN(n660), .Q(n4430), 
        .QN(n1781) );
  DFFR_X1 REGISTERS_reg_2__14_ ( .D(n3512), .CK(CLK), .RN(n660), .Q(n4429), 
        .QN(n1806) );
  DFFR_X1 REGISTERS_reg_2__13_ ( .D(n3511), .CK(CLK), .RN(n660), .Q(n4428), 
        .QN(n1831) );
  DFFR_X1 REGISTERS_reg_2__12_ ( .D(n3510), .CK(CLK), .RN(n659), .Q(n4427), 
        .QN(n1856) );
  DFFR_X1 REGISTERS_reg_2__11_ ( .D(n3509), .CK(CLK), .RN(n659), .Q(n4426), 
        .QN(n1881) );
  DFFR_X1 REGISTERS_reg_2__10_ ( .D(n3508), .CK(CLK), .RN(n659), .Q(n4425), 
        .QN(n1906) );
  DFFR_X1 REGISTERS_reg_2__9_ ( .D(n3507), .CK(CLK), .RN(n659), .Q(n4424), 
        .QN(n1931) );
  DFFR_X1 REGISTERS_reg_2__8_ ( .D(n3506), .CK(CLK), .RN(n659), .Q(n4423), 
        .QN(n1956) );
  DFFR_X1 REGISTERS_reg_2__7_ ( .D(n3505), .CK(CLK), .RN(n659), .Q(n4422), 
        .QN(n1981) );
  DFFR_X1 REGISTERS_reg_2__6_ ( .D(n3504), .CK(CLK), .RN(n659), .Q(n4421), 
        .QN(n2006) );
  DFFR_X1 REGISTERS_reg_2__5_ ( .D(n3503), .CK(CLK), .RN(n659), .Q(n4420), 
        .QN(n2031) );
  DFFR_X1 REGISTERS_reg_2__4_ ( .D(n3502), .CK(CLK), .RN(n659), .Q(n4419), 
        .QN(n2056) );
  DFFR_X1 REGISTERS_reg_2__3_ ( .D(n3501), .CK(CLK), .RN(n659), .Q(n4418), 
        .QN(n2081) );
  DFFR_X1 REGISTERS_reg_2__2_ ( .D(n3500), .CK(CLK), .RN(n659), .Q(n4417), 
        .QN(n2106) );
  DFFR_X1 REGISTERS_reg_2__1_ ( .D(n3499), .CK(CLK), .RN(n659), .Q(n4416), 
        .QN(n2131) );
  DFFR_X1 REGISTERS_reg_2__0_ ( .D(n3498), .CK(CLK), .RN(n658), .Q(n4415), 
        .QN(n2171) );
  DFFR_X1 REGISTERS_reg_15__23_ ( .D(n3105), .CK(CLK), .RN(n646), .Q(n4214) );
  DFFR_X1 REGISTERS_reg_15__22_ ( .D(n3104), .CK(CLK), .RN(n646), .Q(n4213) );
  DFFR_X1 REGISTERS_reg_15__21_ ( .D(n3103), .CK(CLK), .RN(n646), .Q(n4212) );
  DFFR_X1 REGISTERS_reg_15__20_ ( .D(n3102), .CK(CLK), .RN(n646), .Q(n4211) );
  DFFR_X1 REGISTERS_reg_15__19_ ( .D(n3101), .CK(CLK), .RN(n646), .Q(n4210) );
  DFFR_X1 REGISTERS_reg_15__18_ ( .D(n3100), .CK(CLK), .RN(n646), .Q(n4209) );
  DFFR_X1 REGISTERS_reg_15__17_ ( .D(n3099), .CK(CLK), .RN(n646), .Q(n4208) );
  DFFR_X1 REGISTERS_reg_15__16_ ( .D(n3098), .CK(CLK), .RN(n646), .Q(n4207) );
  DFFR_X1 REGISTERS_reg_15__15_ ( .D(n3097), .CK(CLK), .RN(n645), .Q(n4206) );
  DFFR_X1 REGISTERS_reg_15__14_ ( .D(n3096), .CK(CLK), .RN(n645), .Q(n4205) );
  DFFR_X1 REGISTERS_reg_15__13_ ( .D(n3095), .CK(CLK), .RN(n645), .Q(n4204) );
  DFFR_X1 REGISTERS_reg_15__12_ ( .D(n3094), .CK(CLK), .RN(n645), .Q(n4203) );
  DFFR_X1 REGISTERS_reg_15__11_ ( .D(n3093), .CK(CLK), .RN(n645), .Q(n4202) );
  DFFR_X1 REGISTERS_reg_15__10_ ( .D(n3092), .CK(CLK), .RN(n645), .Q(n4201) );
  DFFR_X1 REGISTERS_reg_15__9_ ( .D(n3091), .CK(CLK), .RN(n645), .Q(n4200) );
  DFFR_X1 REGISTERS_reg_15__8_ ( .D(n3090), .CK(CLK), .RN(n645), .Q(n4199) );
  DFFR_X1 REGISTERS_reg_15__7_ ( .D(n3089), .CK(CLK), .RN(n645), .Q(n4198) );
  DFFR_X1 REGISTERS_reg_15__6_ ( .D(n3088), .CK(CLK), .RN(n645), .Q(n4197) );
  DFFR_X1 REGISTERS_reg_15__5_ ( .D(n3087), .CK(CLK), .RN(n645), .Q(n4196) );
  DFFR_X1 REGISTERS_reg_15__4_ ( .D(n3086), .CK(CLK), .RN(n645), .Q(n4195) );
  DFFR_X1 REGISTERS_reg_15__3_ ( .D(n3085), .CK(CLK), .RN(n612), .Q(n4194) );
  DFFR_X1 REGISTERS_reg_15__2_ ( .D(n3084), .CK(CLK), .RN(n612), .Q(n4193) );
  DFFR_X1 REGISTERS_reg_15__1_ ( .D(n3083), .CK(CLK), .RN(n612), .Q(n4192) );
  DFFR_X1 REGISTERS_reg_15__0_ ( .D(n3082), .CK(CLK), .RN(n612), .Q(n4191) );
  DFFR_X1 REGISTERS_reg_14__23_ ( .D(n3137), .CK(CLK), .RN(n649), .Q(n4246) );
  DFFR_X1 REGISTERS_reg_14__22_ ( .D(n3136), .CK(CLK), .RN(n649), .Q(n4245) );
  DFFR_X1 REGISTERS_reg_14__21_ ( .D(n3135), .CK(CLK), .RN(n649), .Q(n4244) );
  DFFR_X1 REGISTERS_reg_14__20_ ( .D(n3134), .CK(CLK), .RN(n649), .Q(n4243) );
  DFFR_X1 REGISTERS_reg_14__19_ ( .D(n3133), .CK(CLK), .RN(n649), .Q(n4242) );
  DFFR_X1 REGISTERS_reg_14__18_ ( .D(n3132), .CK(CLK), .RN(n648), .Q(n4241) );
  DFFR_X1 REGISTERS_reg_14__17_ ( .D(n3131), .CK(CLK), .RN(n648), .Q(n4240) );
  DFFR_X1 REGISTERS_reg_14__16_ ( .D(n3130), .CK(CLK), .RN(n648), .Q(n4239) );
  DFFR_X1 REGISTERS_reg_14__15_ ( .D(n3129), .CK(CLK), .RN(n648), .Q(n4238) );
  DFFR_X1 REGISTERS_reg_14__14_ ( .D(n3128), .CK(CLK), .RN(n648), .Q(n4237) );
  DFFR_X1 REGISTERS_reg_14__13_ ( .D(n3127), .CK(CLK), .RN(n648), .Q(n4236) );
  DFFR_X1 REGISTERS_reg_14__12_ ( .D(n3126), .CK(CLK), .RN(n648), .Q(n4235) );
  DFFR_X1 REGISTERS_reg_14__11_ ( .D(n3125), .CK(CLK), .RN(n648), .Q(n4234) );
  DFFR_X1 REGISTERS_reg_14__10_ ( .D(n3124), .CK(CLK), .RN(n648), .Q(n4233) );
  DFFR_X1 REGISTERS_reg_14__9_ ( .D(n3123), .CK(CLK), .RN(n648), .Q(n4232) );
  DFFR_X1 REGISTERS_reg_14__8_ ( .D(n3122), .CK(CLK), .RN(n648), .Q(n4231) );
  DFFR_X1 REGISTERS_reg_14__7_ ( .D(n3121), .CK(CLK), .RN(n647), .Q(n4230) );
  DFFR_X1 REGISTERS_reg_14__6_ ( .D(n3120), .CK(CLK), .RN(n647), .Q(n4229) );
  DFFR_X1 REGISTERS_reg_14__5_ ( .D(n3119), .CK(CLK), .RN(n647), .Q(n4228) );
  DFFR_X1 REGISTERS_reg_14__4_ ( .D(n3118), .CK(CLK), .RN(n647), .Q(n4227) );
  DFFR_X1 REGISTERS_reg_14__3_ ( .D(n3117), .CK(CLK), .RN(n647), .Q(n4226) );
  DFFR_X1 REGISTERS_reg_14__2_ ( .D(n3116), .CK(CLK), .RN(n647), .Q(n4225) );
  DFFR_X1 REGISTERS_reg_14__1_ ( .D(n3115), .CK(CLK), .RN(n647), .Q(n4224) );
  DFFR_X1 REGISTERS_reg_14__0_ ( .D(n3114), .CK(CLK), .RN(n647), .Q(n4223) );
  DFFR_X1 REGISTERS_reg_23__23_ ( .D(n2849), .CK(CLK), .RN(n707), .Q(n4086), 
        .QN(n1563) );
  DFFR_X1 REGISTERS_reg_23__22_ ( .D(n2848), .CK(CLK), .RN(n707), .Q(n4085), 
        .QN(n1588) );
  DFFR_X1 REGISTERS_reg_23__21_ ( .D(n2847), .CK(CLK), .RN(n707), .Q(n4084), 
        .QN(n1613) );
  DFFR_X1 REGISTERS_reg_23__20_ ( .D(n2846), .CK(CLK), .RN(n707), .Q(n4083), 
        .QN(n1638) );
  DFFR_X1 REGISTERS_reg_23__19_ ( .D(n2845), .CK(CLK), .RN(n707), .Q(n4082), 
        .QN(n1663) );
  DFFR_X1 REGISTERS_reg_23__18_ ( .D(n2844), .CK(CLK), .RN(n707), .Q(n4081), 
        .QN(n1688) );
  DFFR_X1 REGISTERS_reg_23__17_ ( .D(n2843), .CK(CLK), .RN(n707), .Q(n4080), 
        .QN(n1713) );
  DFFR_X1 REGISTERS_reg_23__16_ ( .D(n2842), .CK(CLK), .RN(n707), .Q(n4079), 
        .QN(n1738) );
  DFFR_X1 REGISTERS_reg_23__15_ ( .D(n2841), .CK(CLK), .RN(n707), .Q(n4078), 
        .QN(n1763) );
  DFFR_X1 REGISTERS_reg_23__14_ ( .D(n2840), .CK(CLK), .RN(n707), .Q(n4077), 
        .QN(n1788) );
  DFFR_X1 REGISTERS_reg_23__13_ ( .D(n2839), .CK(CLK), .RN(n707), .Q(n4076), 
        .QN(n1813) );
  DFFR_X1 REGISTERS_reg_23__12_ ( .D(n2838), .CK(CLK), .RN(n707), .Q(n4075), 
        .QN(n1838) );
  DFFR_X1 REGISTERS_reg_23__11_ ( .D(n2837), .CK(CLK), .RN(n706), .Q(n4074), 
        .QN(n1863) );
  DFFR_X1 REGISTERS_reg_23__10_ ( .D(n2836), .CK(CLK), .RN(n706), .Q(n4073), 
        .QN(n1888) );
  DFFR_X1 REGISTERS_reg_23__9_ ( .D(n2835), .CK(CLK), .RN(n706), .Q(n4072), 
        .QN(n1913) );
  DFFR_X1 REGISTERS_reg_23__8_ ( .D(n2834), .CK(CLK), .RN(n706), .Q(n4071), 
        .QN(n1938) );
  DFFR_X1 REGISTERS_reg_23__7_ ( .D(n2833), .CK(CLK), .RN(n706), .Q(n4070), 
        .QN(n1963) );
  DFFR_X1 REGISTERS_reg_23__6_ ( .D(n2832), .CK(CLK), .RN(n706), .Q(n4069), 
        .QN(n1988) );
  DFFR_X1 REGISTERS_reg_23__5_ ( .D(n2831), .CK(CLK), .RN(n706), .Q(n4068), 
        .QN(n2013) );
  DFFR_X1 REGISTERS_reg_23__4_ ( .D(n2830), .CK(CLK), .RN(n706), .Q(n4067), 
        .QN(n2038) );
  DFFR_X1 REGISTERS_reg_23__3_ ( .D(n2829), .CK(CLK), .RN(n706), .Q(n4066), 
        .QN(n2063) );
  DFFR_X1 REGISTERS_reg_23__2_ ( .D(n2828), .CK(CLK), .RN(n706), .Q(n4065), 
        .QN(n2088) );
  DFFR_X1 REGISTERS_reg_23__1_ ( .D(n2827), .CK(CLK), .RN(n706), .Q(n4064), 
        .QN(n2113) );
  DFFR_X1 REGISTERS_reg_23__0_ ( .D(n2826), .CK(CLK), .RN(n706), .Q(n4063), 
        .QN(n2139) );
  DFFR_X1 REGISTERS_reg_22__23_ ( .D(n2881), .CK(CLK), .RN(n710), .Q(n4118), 
        .QN(n1570) );
  DFFR_X1 REGISTERS_reg_22__22_ ( .D(n2880), .CK(CLK), .RN(n710), .Q(n4117), 
        .QN(n1595) );
  DFFR_X1 REGISTERS_reg_22__21_ ( .D(n2879), .CK(CLK), .RN(n710), .Q(n4116), 
        .QN(n1620) );
  DFFR_X1 REGISTERS_reg_22__20_ ( .D(n2878), .CK(CLK), .RN(n710), .Q(n4115), 
        .QN(n1645) );
  DFFR_X1 REGISTERS_reg_22__19_ ( .D(n2877), .CK(CLK), .RN(n710), .Q(n4114), 
        .QN(n1670) );
  DFFR_X1 REGISTERS_reg_22__18_ ( .D(n2876), .CK(CLK), .RN(n710), .Q(n4113), 
        .QN(n1695) );
  DFFR_X1 REGISTERS_reg_22__17_ ( .D(n2875), .CK(CLK), .RN(n710), .Q(n4112), 
        .QN(n1720) );
  DFFR_X1 REGISTERS_reg_22__16_ ( .D(n2874), .CK(CLK), .RN(n710), .Q(n4111), 
        .QN(n1745) );
  DFFR_X1 REGISTERS_reg_22__15_ ( .D(n2873), .CK(CLK), .RN(n709), .Q(n4110), 
        .QN(n1770) );
  DFFR_X1 REGISTERS_reg_22__14_ ( .D(n2872), .CK(CLK), .RN(n709), .Q(n4109), 
        .QN(n1795) );
  DFFR_X1 REGISTERS_reg_22__13_ ( .D(n2871), .CK(CLK), .RN(n709), .Q(n4108), 
        .QN(n1820) );
  DFFR_X1 REGISTERS_reg_22__12_ ( .D(n2870), .CK(CLK), .RN(n709), .Q(n4107), 
        .QN(n1845) );
  DFFR_X1 REGISTERS_reg_22__11_ ( .D(n2869), .CK(CLK), .RN(n709), .Q(n4106), 
        .QN(n1870) );
  DFFR_X1 REGISTERS_reg_22__10_ ( .D(n2868), .CK(CLK), .RN(n709), .Q(n4105), 
        .QN(n1895) );
  DFFR_X1 REGISTERS_reg_22__9_ ( .D(n2867), .CK(CLK), .RN(n709), .Q(n4104), 
        .QN(n1920) );
  DFFR_X1 REGISTERS_reg_22__8_ ( .D(n2866), .CK(CLK), .RN(n709), .Q(n4103), 
        .QN(n1945) );
  DFFR_X1 REGISTERS_reg_22__7_ ( .D(n2865), .CK(CLK), .RN(n709), .Q(n4102), 
        .QN(n1970) );
  DFFR_X1 REGISTERS_reg_22__6_ ( .D(n2864), .CK(CLK), .RN(n709), .Q(n4101), 
        .QN(n1995) );
  DFFR_X1 REGISTERS_reg_22__5_ ( .D(n2863), .CK(CLK), .RN(n709), .Q(n4100), 
        .QN(n2020) );
  DFFR_X1 REGISTERS_reg_22__4_ ( .D(n2862), .CK(CLK), .RN(n709), .Q(n4099), 
        .QN(n2045) );
  DFFR_X1 REGISTERS_reg_22__3_ ( .D(n2861), .CK(CLK), .RN(n708), .Q(n4098), 
        .QN(n2070) );
  DFFR_X1 REGISTERS_reg_22__2_ ( .D(n2860), .CK(CLK), .RN(n708), .Q(n4097), 
        .QN(n2095) );
  DFFR_X1 REGISTERS_reg_22__1_ ( .D(n2859), .CK(CLK), .RN(n708), .Q(n4096), 
        .QN(n2120) );
  DFFR_X1 REGISTERS_reg_22__0_ ( .D(n2858), .CK(CLK), .RN(n708), .Q(n4095), 
        .QN(n2155) );
  DFFR_X1 REGISTERS_reg_11__23_ ( .D(n3233), .CK(CLK), .RN(n604), .Q(n4278) );
  DFFR_X1 REGISTERS_reg_11__22_ ( .D(n3232), .CK(CLK), .RN(n604), .Q(n4277) );
  DFFR_X1 REGISTERS_reg_11__21_ ( .D(n3231), .CK(CLK), .RN(n604), .Q(n4276) );
  DFFR_X1 REGISTERS_reg_11__20_ ( .D(n3230), .CK(CLK), .RN(n604), .Q(n4275) );
  DFFR_X1 REGISTERS_reg_11__19_ ( .D(n3229), .CK(CLK), .RN(n604), .Q(n4274) );
  DFFR_X1 REGISTERS_reg_11__18_ ( .D(n3228), .CK(CLK), .RN(n604), .Q(n4273) );
  DFFR_X1 REGISTERS_reg_11__17_ ( .D(n3227), .CK(CLK), .RN(n604), .Q(n4272) );
  DFFR_X1 REGISTERS_reg_11__16_ ( .D(n3226), .CK(CLK), .RN(n604), .Q(n4271) );
  DFFR_X1 REGISTERS_reg_11__15_ ( .D(n3225), .CK(CLK), .RN(n604), .Q(n4270) );
  DFFR_X1 REGISTERS_reg_11__14_ ( .D(n3224), .CK(CLK), .RN(n603), .Q(n4269) );
  DFFR_X1 REGISTERS_reg_11__13_ ( .D(n3223), .CK(CLK), .RN(n603), .Q(n4268) );
  DFFR_X1 REGISTERS_reg_11__12_ ( .D(n3222), .CK(CLK), .RN(n603), .Q(n4267) );
  DFFR_X1 REGISTERS_reg_11__11_ ( .D(n3221), .CK(CLK), .RN(n603), .Q(n4266) );
  DFFR_X1 REGISTERS_reg_11__10_ ( .D(n3220), .CK(CLK), .RN(n603), .Q(n4265) );
  DFFR_X1 REGISTERS_reg_11__9_ ( .D(n3219), .CK(CLK), .RN(n603), .Q(n4264) );
  DFFR_X1 REGISTERS_reg_11__8_ ( .D(n3218), .CK(CLK), .RN(n603), .Q(n4263) );
  DFFR_X1 REGISTERS_reg_11__7_ ( .D(n3217), .CK(CLK), .RN(n603), .Q(n4262) );
  DFFR_X1 REGISTERS_reg_11__6_ ( .D(n3216), .CK(CLK), .RN(n603), .Q(n4261) );
  DFFR_X1 REGISTERS_reg_11__5_ ( .D(n3215), .CK(CLK), .RN(n603), .Q(n4260) );
  DFFR_X1 REGISTERS_reg_11__4_ ( .D(n3214), .CK(CLK), .RN(n603), .Q(n4259) );
  DFFR_X1 REGISTERS_reg_11__3_ ( .D(n3213), .CK(CLK), .RN(n603), .Q(n4258) );
  DFFR_X1 REGISTERS_reg_11__2_ ( .D(n3212), .CK(CLK), .RN(n602), .Q(n4257) );
  DFFR_X1 REGISTERS_reg_11__1_ ( .D(n3211), .CK(CLK), .RN(n602), .Q(n4256) );
  DFFR_X1 REGISTERS_reg_11__0_ ( .D(n3210), .CK(CLK), .RN(n602), .Q(n4255) );
  DFFR_X1 REGISTERS_reg_10__23_ ( .D(n3265), .CK(CLK), .RN(n607), .Q(n4310) );
  DFFR_X1 REGISTERS_reg_10__22_ ( .D(n3264), .CK(CLK), .RN(n607), .Q(n4309) );
  DFFR_X1 REGISTERS_reg_10__21_ ( .D(n3263), .CK(CLK), .RN(n607), .Q(n4308) );
  DFFR_X1 REGISTERS_reg_10__20_ ( .D(n3262), .CK(CLK), .RN(n607), .Q(n4307) );
  DFFR_X1 REGISTERS_reg_10__19_ ( .D(n3261), .CK(CLK), .RN(n607), .Q(n4306) );
  DFFR_X1 REGISTERS_reg_10__18_ ( .D(n3260), .CK(CLK), .RN(n607), .Q(n4305) );
  DFFR_X1 REGISTERS_reg_10__17_ ( .D(n3259), .CK(CLK), .RN(n606), .Q(n4304) );
  DFFR_X1 REGISTERS_reg_10__16_ ( .D(n3258), .CK(CLK), .RN(n606), .Q(n4303) );
  DFFR_X1 REGISTERS_reg_10__15_ ( .D(n3257), .CK(CLK), .RN(n606), .Q(n4302) );
  DFFR_X1 REGISTERS_reg_10__14_ ( .D(n3256), .CK(CLK), .RN(n606), .Q(n4301) );
  DFFR_X1 REGISTERS_reg_10__13_ ( .D(n3255), .CK(CLK), .RN(n606), .Q(n4300) );
  DFFR_X1 REGISTERS_reg_10__12_ ( .D(n3254), .CK(CLK), .RN(n606), .Q(n4299) );
  DFFR_X1 REGISTERS_reg_10__11_ ( .D(n3253), .CK(CLK), .RN(n606), .Q(n4298) );
  DFFR_X1 REGISTERS_reg_10__10_ ( .D(n3252), .CK(CLK), .RN(n606), .Q(n4297) );
  DFFR_X1 REGISTERS_reg_10__9_ ( .D(n3251), .CK(CLK), .RN(n606), .Q(n4296) );
  DFFR_X1 REGISTERS_reg_10__8_ ( .D(n3250), .CK(CLK), .RN(n606), .Q(n4295) );
  DFFR_X1 REGISTERS_reg_10__7_ ( .D(n3249), .CK(CLK), .RN(n606), .Q(n4294) );
  DFFR_X1 REGISTERS_reg_10__6_ ( .D(n3248), .CK(CLK), .RN(n605), .Q(n4293) );
  DFFR_X1 REGISTERS_reg_10__5_ ( .D(n3247), .CK(CLK), .RN(n605), .Q(n4292) );
  DFFR_X1 REGISTERS_reg_10__4_ ( .D(n3246), .CK(CLK), .RN(n605), .Q(n4291) );
  DFFR_X1 REGISTERS_reg_10__3_ ( .D(n3245), .CK(CLK), .RN(n605), .Q(n4290) );
  DFFR_X1 REGISTERS_reg_10__2_ ( .D(n3244), .CK(CLK), .RN(n605), .Q(n4289) );
  DFFR_X1 REGISTERS_reg_10__1_ ( .D(n3243), .CK(CLK), .RN(n605), .Q(n4288) );
  DFFR_X1 REGISTERS_reg_10__0_ ( .D(n3242), .CK(CLK), .RN(n605), .Q(n4287) );
  DFFR_X1 REGISTERS_reg_19__23_ ( .D(n2977), .CK(CLK), .RN(n698), .Q(n4150) );
  DFFR_X1 REGISTERS_reg_19__22_ ( .D(n2976), .CK(CLK), .RN(n697), .Q(n4149) );
  DFFR_X1 REGISTERS_reg_19__21_ ( .D(n2975), .CK(CLK), .RN(n697), .Q(n4148) );
  DFFR_X1 REGISTERS_reg_19__20_ ( .D(n2974), .CK(CLK), .RN(n697), .Q(n4147) );
  DFFR_X1 REGISTERS_reg_19__19_ ( .D(n2973), .CK(CLK), .RN(n697), .Q(n4146) );
  DFFR_X1 REGISTERS_reg_19__18_ ( .D(n2972), .CK(CLK), .RN(n697), .Q(n4145) );
  DFFR_X1 REGISTERS_reg_19__17_ ( .D(n2971), .CK(CLK), .RN(n697), .Q(n4144) );
  DFFR_X1 REGISTERS_reg_19__16_ ( .D(n2970), .CK(CLK), .RN(n697), .Q(n4143) );
  DFFR_X1 REGISTERS_reg_19__15_ ( .D(n2969), .CK(CLK), .RN(n697), .Q(n4142) );
  DFFR_X1 REGISTERS_reg_19__14_ ( .D(n2968), .CK(CLK), .RN(n697), .Q(n4141) );
  DFFR_X1 REGISTERS_reg_19__13_ ( .D(n2967), .CK(CLK), .RN(n697), .Q(n4140) );
  DFFR_X1 REGISTERS_reg_19__12_ ( .D(n2966), .CK(CLK), .RN(n697), .Q(n4139) );
  DFFR_X1 REGISTERS_reg_19__11_ ( .D(n2965), .CK(CLK), .RN(n697), .Q(n4138) );
  DFFR_X1 REGISTERS_reg_19__10_ ( .D(n2964), .CK(CLK), .RN(n696), .Q(n4137) );
  DFFR_X1 REGISTERS_reg_19__9_ ( .D(n2963), .CK(CLK), .RN(n696), .Q(n4136) );
  DFFR_X1 REGISTERS_reg_19__8_ ( .D(n2962), .CK(CLK), .RN(n696), .Q(n4135) );
  DFFR_X1 REGISTERS_reg_19__7_ ( .D(n2961), .CK(CLK), .RN(n696), .Q(n4134) );
  DFFR_X1 REGISTERS_reg_19__6_ ( .D(n2960), .CK(CLK), .RN(n696), .Q(n4133) );
  DFFR_X1 REGISTERS_reg_19__5_ ( .D(n2959), .CK(CLK), .RN(n696), .Q(n4132) );
  DFFR_X1 REGISTERS_reg_19__4_ ( .D(n2958), .CK(CLK), .RN(n696), .Q(n4131) );
  DFFR_X1 REGISTERS_reg_19__3_ ( .D(n2957), .CK(CLK), .RN(n696), .Q(n4130) );
  DFFR_X1 REGISTERS_reg_19__2_ ( .D(n2956), .CK(CLK), .RN(n696), .Q(n4129) );
  DFFR_X1 REGISTERS_reg_19__1_ ( .D(n2955), .CK(CLK), .RN(n696), .Q(n4128) );
  DFFR_X1 REGISTERS_reg_19__0_ ( .D(n2954), .CK(CLK), .RN(n696), .Q(n4127) );
  DFFR_X1 REGISTERS_reg_18__23_ ( .D(n3009), .CK(CLK), .RN(n700), .Q(n4182) );
  DFFR_X1 REGISTERS_reg_18__22_ ( .D(n3008), .CK(CLK), .RN(n700), .Q(n4181) );
  DFFR_X1 REGISTERS_reg_18__21_ ( .D(n3007), .CK(CLK), .RN(n700), .Q(n4180) );
  DFFR_X1 REGISTERS_reg_18__20_ ( .D(n3006), .CK(CLK), .RN(n700), .Q(n4179) );
  DFFR_X1 REGISTERS_reg_18__19_ ( .D(n3005), .CK(CLK), .RN(n700), .Q(n4178) );
  DFFR_X1 REGISTERS_reg_18__18_ ( .D(n3004), .CK(CLK), .RN(n700), .Q(n4177) );
  DFFR_X1 REGISTERS_reg_18__17_ ( .D(n3003), .CK(CLK), .RN(n700), .Q(n4176) );
  DFFR_X1 REGISTERS_reg_18__16_ ( .D(n3002), .CK(CLK), .RN(n700), .Q(n4175) );
  DFFR_X1 REGISTERS_reg_18__15_ ( .D(n3001), .CK(CLK), .RN(n700), .Q(n4174) );
  DFFR_X1 REGISTERS_reg_18__14_ ( .D(n3000), .CK(CLK), .RN(n699), .Q(n4173) );
  DFFR_X1 REGISTERS_reg_18__13_ ( .D(n2999), .CK(CLK), .RN(n699), .Q(n4172) );
  DFFR_X1 REGISTERS_reg_18__12_ ( .D(n2998), .CK(CLK), .RN(n699), .Q(n4171) );
  DFFR_X1 REGISTERS_reg_18__11_ ( .D(n2997), .CK(CLK), .RN(n699), .Q(n4170) );
  DFFR_X1 REGISTERS_reg_18__10_ ( .D(n2996), .CK(CLK), .RN(n699), .Q(n4169) );
  DFFR_X1 REGISTERS_reg_18__9_ ( .D(n2995), .CK(CLK), .RN(n699), .Q(n4168) );
  DFFR_X1 REGISTERS_reg_18__8_ ( .D(n2994), .CK(CLK), .RN(n699), .Q(n4167) );
  DFFR_X1 REGISTERS_reg_18__7_ ( .D(n2993), .CK(CLK), .RN(n699), .Q(n4166) );
  DFFR_X1 REGISTERS_reg_18__6_ ( .D(n2992), .CK(CLK), .RN(n699), .Q(n4165) );
  DFFR_X1 REGISTERS_reg_18__5_ ( .D(n2991), .CK(CLK), .RN(n699), .Q(n4164) );
  DFFR_X1 REGISTERS_reg_18__4_ ( .D(n2990), .CK(CLK), .RN(n699), .Q(n4163) );
  DFFR_X1 REGISTERS_reg_18__3_ ( .D(n2989), .CK(CLK), .RN(n699), .Q(n4162) );
  DFFR_X1 REGISTERS_reg_18__2_ ( .D(n2988), .CK(CLK), .RN(n698), .Q(n4161) );
  DFFR_X1 REGISTERS_reg_18__1_ ( .D(n2987), .CK(CLK), .RN(n698), .Q(n4160) );
  DFFR_X1 REGISTERS_reg_18__0_ ( .D(n2986), .CK(CLK), .RN(n698), .Q(n4159) );
  DFFR_X1 REGISTERS_reg_29__23_ ( .D(n2657), .CK(CLK), .RN(n692), .Q(n3958) );
  DFFR_X1 REGISTERS_reg_29__22_ ( .D(n2656), .CK(CLK), .RN(n691), .Q(n3957) );
  DFFR_X1 REGISTERS_reg_29__21_ ( .D(n2655), .CK(CLK), .RN(n691), .Q(n3956) );
  DFFR_X1 REGISTERS_reg_29__20_ ( .D(n2654), .CK(CLK), .RN(n691), .Q(n3955) );
  DFFR_X1 REGISTERS_reg_29__19_ ( .D(n2653), .CK(CLK), .RN(n691), .Q(n3954) );
  DFFR_X1 REGISTERS_reg_29__18_ ( .D(n2652), .CK(CLK), .RN(n691), .Q(n3953) );
  DFFR_X1 REGISTERS_reg_29__17_ ( .D(n2651), .CK(CLK), .RN(n691), .Q(n3952) );
  DFFR_X1 REGISTERS_reg_29__16_ ( .D(n2650), .CK(CLK), .RN(n691), .Q(n3951) );
  DFFR_X1 REGISTERS_reg_29__15_ ( .D(n2649), .CK(CLK), .RN(n691), .Q(n3950) );
  DFFR_X1 REGISTERS_reg_29__14_ ( .D(n2648), .CK(CLK), .RN(n691), .Q(n3949) );
  DFFR_X1 REGISTERS_reg_29__13_ ( .D(n2647), .CK(CLK), .RN(n691), .Q(n3948) );
  DFFR_X1 REGISTERS_reg_29__12_ ( .D(n2646), .CK(CLK), .RN(n691), .Q(n3947) );
  DFFR_X1 REGISTERS_reg_29__11_ ( .D(n2645), .CK(CLK), .RN(n691), .Q(n3946) );
  DFFR_X1 REGISTERS_reg_29__10_ ( .D(n2644), .CK(CLK), .RN(n690), .Q(n3945) );
  DFFR_X1 REGISTERS_reg_29__9_ ( .D(n2643), .CK(CLK), .RN(n690), .Q(n3944) );
  DFFR_X1 REGISTERS_reg_29__8_ ( .D(n2642), .CK(CLK), .RN(n690), .Q(n3943) );
  DFFR_X1 REGISTERS_reg_29__7_ ( .D(n2641), .CK(CLK), .RN(n690), .Q(n3942) );
  DFFR_X1 REGISTERS_reg_29__6_ ( .D(n2640), .CK(CLK), .RN(n690), .Q(n3941) );
  DFFR_X1 REGISTERS_reg_29__5_ ( .D(n2639), .CK(CLK), .RN(n690), .Q(n3940) );
  DFFR_X1 REGISTERS_reg_29__4_ ( .D(n2638), .CK(CLK), .RN(n690), .Q(n3939) );
  DFFR_X1 REGISTERS_reg_29__3_ ( .D(n2637), .CK(CLK), .RN(n690), .Q(n3938) );
  DFFR_X1 REGISTERS_reg_29__2_ ( .D(n2636), .CK(CLK), .RN(n690), .Q(n3937) );
  DFFR_X1 REGISTERS_reg_29__1_ ( .D(n2635), .CK(CLK), .RN(n690), .Q(n3936) );
  DFFR_X1 REGISTERS_reg_29__0_ ( .D(n2634), .CK(CLK), .RN(n690), .Q(n3935) );
  DFFR_X1 REGISTERS_reg_28__23_ ( .D(n2689), .CK(CLK), .RN(n694), .Q(n3990), 
        .QN(n1565) );
  DFFR_X1 REGISTERS_reg_28__22_ ( .D(n2688), .CK(CLK), .RN(n694), .Q(n3989), 
        .QN(n1590) );
  DFFR_X1 REGISTERS_reg_28__21_ ( .D(n2687), .CK(CLK), .RN(n694), .Q(n3988), 
        .QN(n1615) );
  DFFR_X1 REGISTERS_reg_28__20_ ( .D(n2686), .CK(CLK), .RN(n694), .Q(n3987), 
        .QN(n1640) );
  DFFR_X1 REGISTERS_reg_28__19_ ( .D(n2685), .CK(CLK), .RN(n694), .Q(n3986), 
        .QN(n1665) );
  DFFR_X1 REGISTERS_reg_28__18_ ( .D(n2684), .CK(CLK), .RN(n694), .Q(n3985), 
        .QN(n1690) );
  DFFR_X1 REGISTERS_reg_28__17_ ( .D(n2683), .CK(CLK), .RN(n694), .Q(n3984), 
        .QN(n1715) );
  DFFR_X1 REGISTERS_reg_28__16_ ( .D(n2682), .CK(CLK), .RN(n694), .Q(n3983), 
        .QN(n1740) );
  DFFR_X1 REGISTERS_reg_28__15_ ( .D(n2681), .CK(CLK), .RN(n694), .Q(n3982), 
        .QN(n1765) );
  DFFR_X1 REGISTERS_reg_28__14_ ( .D(n2680), .CK(CLK), .RN(n693), .Q(n3981), 
        .QN(n1790) );
  DFFR_X1 REGISTERS_reg_28__13_ ( .D(n2679), .CK(CLK), .RN(n693), .Q(n3980), 
        .QN(n1815) );
  DFFR_X1 REGISTERS_reg_28__12_ ( .D(n2678), .CK(CLK), .RN(n693), .Q(n3979), 
        .QN(n1840) );
  DFFR_X1 REGISTERS_reg_28__11_ ( .D(n2677), .CK(CLK), .RN(n693), .Q(n3978), 
        .QN(n1865) );
  DFFR_X1 REGISTERS_reg_28__10_ ( .D(n2676), .CK(CLK), .RN(n693), .Q(n3977), 
        .QN(n1890) );
  DFFR_X1 REGISTERS_reg_28__9_ ( .D(n2675), .CK(CLK), .RN(n693), .Q(n3976), 
        .QN(n1915) );
  DFFR_X1 REGISTERS_reg_28__8_ ( .D(n2674), .CK(CLK), .RN(n693), .Q(n3975), 
        .QN(n1940) );
  DFFR_X1 REGISTERS_reg_28__7_ ( .D(n2673), .CK(CLK), .RN(n693), .Q(n3974), 
        .QN(n1965) );
  DFFR_X1 REGISTERS_reg_28__6_ ( .D(n2672), .CK(CLK), .RN(n693), .Q(n3973), 
        .QN(n1990) );
  DFFR_X1 REGISTERS_reg_28__5_ ( .D(n2671), .CK(CLK), .RN(n693), .Q(n3972), 
        .QN(n2015) );
  DFFR_X1 REGISTERS_reg_28__4_ ( .D(n2670), .CK(CLK), .RN(n693), .Q(n3971), 
        .QN(n2040) );
  DFFR_X1 REGISTERS_reg_28__3_ ( .D(n2669), .CK(CLK), .RN(n693), .Q(n3970), 
        .QN(n2065) );
  DFFR_X1 REGISTERS_reg_28__2_ ( .D(n2668), .CK(CLK), .RN(n692), .Q(n3969), 
        .QN(n2090) );
  DFFR_X1 REGISTERS_reg_28__1_ ( .D(n2667), .CK(CLK), .RN(n692), .Q(n3968), 
        .QN(n2115) );
  DFFR_X1 REGISTERS_reg_28__0_ ( .D(n2666), .CK(CLK), .RN(n692), .Q(n3967), 
        .QN(n2147) );
  DFFR_X1 REGISTERS_reg_25__23_ ( .D(n2785), .CK(CLK), .RN(n682), .Q(n4022) );
  DFFR_X1 REGISTERS_reg_25__22_ ( .D(n2784), .CK(CLK), .RN(n681), .Q(n4021) );
  DFFR_X1 REGISTERS_reg_25__21_ ( .D(n2783), .CK(CLK), .RN(n681), .Q(n4020) );
  DFFR_X1 REGISTERS_reg_25__20_ ( .D(n2782), .CK(CLK), .RN(n681), .Q(n4019) );
  DFFR_X1 REGISTERS_reg_25__19_ ( .D(n2781), .CK(CLK), .RN(n681), .Q(n4018) );
  DFFR_X1 REGISTERS_reg_25__18_ ( .D(n2780), .CK(CLK), .RN(n681), .Q(n4017) );
  DFFR_X1 REGISTERS_reg_25__17_ ( .D(n2779), .CK(CLK), .RN(n681), .Q(n4016) );
  DFFR_X1 REGISTERS_reg_25__16_ ( .D(n2778), .CK(CLK), .RN(n681), .Q(n4015) );
  DFFR_X1 REGISTERS_reg_25__15_ ( .D(n2777), .CK(CLK), .RN(n681), .Q(n4014) );
  DFFR_X1 REGISTERS_reg_25__14_ ( .D(n2776), .CK(CLK), .RN(n681), .Q(n4013) );
  DFFR_X1 REGISTERS_reg_25__13_ ( .D(n2775), .CK(CLK), .RN(n681), .Q(n4012) );
  DFFR_X1 REGISTERS_reg_25__12_ ( .D(n2774), .CK(CLK), .RN(n681), .Q(n4011) );
  DFFR_X1 REGISTERS_reg_25__11_ ( .D(n2773), .CK(CLK), .RN(n681), .Q(n4010) );
  DFFR_X1 REGISTERS_reg_25__10_ ( .D(n2772), .CK(CLK), .RN(n680), .Q(n4009) );
  DFFR_X1 REGISTERS_reg_25__9_ ( .D(n2771), .CK(CLK), .RN(n680), .Q(n4008) );
  DFFR_X1 REGISTERS_reg_25__8_ ( .D(n2770), .CK(CLK), .RN(n680), .Q(n4007) );
  DFFR_X1 REGISTERS_reg_25__7_ ( .D(n2769), .CK(CLK), .RN(n680), .Q(n4006) );
  DFFR_X1 REGISTERS_reg_25__6_ ( .D(n2768), .CK(CLK), .RN(n680), .Q(n4005) );
  DFFR_X1 REGISTERS_reg_25__5_ ( .D(n2767), .CK(CLK), .RN(n680), .Q(n4004) );
  DFFR_X1 REGISTERS_reg_25__4_ ( .D(n2766), .CK(CLK), .RN(n680), .Q(n4003) );
  DFFR_X1 REGISTERS_reg_25__3_ ( .D(n2765), .CK(CLK), .RN(n680), .Q(n4002) );
  DFFR_X1 REGISTERS_reg_25__2_ ( .D(n2764), .CK(CLK), .RN(n680), .Q(n4001) );
  DFFR_X1 REGISTERS_reg_25__1_ ( .D(n2763), .CK(CLK), .RN(n680), .Q(n4000) );
  DFFR_X1 REGISTERS_reg_25__0_ ( .D(n2762), .CK(CLK), .RN(n680), .Q(n3999) );
  DFFR_X1 REGISTERS_reg_24__23_ ( .D(n2817), .CK(CLK), .RN(n684), .Q(n4054) );
  DFFR_X1 REGISTERS_reg_24__22_ ( .D(n2816), .CK(CLK), .RN(n684), .Q(n4053) );
  DFFR_X1 REGISTERS_reg_24__21_ ( .D(n2815), .CK(CLK), .RN(n684), .Q(n4052) );
  DFFR_X1 REGISTERS_reg_24__20_ ( .D(n2814), .CK(CLK), .RN(n684), .Q(n4051) );
  DFFR_X1 REGISTERS_reg_24__19_ ( .D(n2813), .CK(CLK), .RN(n684), .Q(n4050) );
  DFFR_X1 REGISTERS_reg_24__18_ ( .D(n2812), .CK(CLK), .RN(n684), .Q(n4049) );
  DFFR_X1 REGISTERS_reg_24__17_ ( .D(n2811), .CK(CLK), .RN(n684), .Q(n4048) );
  DFFR_X1 REGISTERS_reg_24__16_ ( .D(n2810), .CK(CLK), .RN(n684), .Q(n4047) );
  DFFR_X1 REGISTERS_reg_24__15_ ( .D(n2809), .CK(CLK), .RN(n684), .Q(n4046) );
  DFFR_X1 REGISTERS_reg_24__14_ ( .D(n2808), .CK(CLK), .RN(n683), .Q(n4045) );
  DFFR_X1 REGISTERS_reg_24__13_ ( .D(n2807), .CK(CLK), .RN(n683), .Q(n4044) );
  DFFR_X1 REGISTERS_reg_24__12_ ( .D(n2806), .CK(CLK), .RN(n683), .Q(n4043) );
  DFFR_X1 REGISTERS_reg_24__11_ ( .D(n2805), .CK(CLK), .RN(n683), .Q(n4042) );
  DFFR_X1 REGISTERS_reg_24__10_ ( .D(n2804), .CK(CLK), .RN(n683), .Q(n4041) );
  DFFR_X1 REGISTERS_reg_24__9_ ( .D(n2803), .CK(CLK), .RN(n683), .Q(n4040) );
  DFFR_X1 REGISTERS_reg_24__8_ ( .D(n2802), .CK(CLK), .RN(n683), .Q(n4039) );
  DFFR_X1 REGISTERS_reg_24__7_ ( .D(n2801), .CK(CLK), .RN(n683), .Q(n4038) );
  DFFR_X1 REGISTERS_reg_24__6_ ( .D(n2800), .CK(CLK), .RN(n683), .Q(n4037) );
  DFFR_X1 REGISTERS_reg_24__5_ ( .D(n2799), .CK(CLK), .RN(n683), .Q(n4036) );
  DFFR_X1 REGISTERS_reg_24__4_ ( .D(n2798), .CK(CLK), .RN(n683), .Q(n4035) );
  DFF_X1 OUT1_reg_8_ ( .D(n2514), .CK(CLK), .Q(OUT1[8]), .QN(n3879) );
  DFF_X1 OUT1_reg_2_ ( .D(n2508), .CK(CLK), .Q(OUT1[2]), .QN(n3873) );
  DFF_X1 OUT1_reg_13_ ( .D(n2519), .CK(CLK), .Q(OUT1[13]), .QN(n3884) );
  DFF_X1 OUT1_reg_12_ ( .D(n2518), .CK(CLK), .Q(OUT1[12]), .QN(n3883) );
  DFF_X1 OUT1_reg_9_ ( .D(n2515), .CK(CLK), .Q(OUT1[9]), .QN(n3880) );
  DFF_X1 OUT1_reg_4_ ( .D(n2510), .CK(CLK), .Q(OUT1[4]), .QN(n3875) );
  DFF_X1 OUT1_reg_3_ ( .D(n2509), .CK(CLK), .Q(OUT1[3]), .QN(n3874) );
  DFF_X1 OUT1_reg_1_ ( .D(n2507), .CK(CLK), .Q(OUT1[1]), .QN(n3872) );
  DFF_X1 OUT1_reg_17_ ( .D(n2523), .CK(CLK), .Q(OUT1[17]), .QN(n3888) );
  DFF_X1 OUT1_reg_16_ ( .D(n2522), .CK(CLK), .Q(OUT1[16]), .QN(n3887) );
  DFF_X1 OUT1_reg_15_ ( .D(n2521), .CK(CLK), .Q(OUT1[15]), .QN(n3886) );
  DFF_X1 OUT1_reg_14_ ( .D(n2520), .CK(CLK), .Q(OUT1[14]), .QN(n3885) );
  DFF_X1 OUT2_reg_10_ ( .D(n2548), .CK(CLK), .Q(OUT2[10]), .QN(n3913) );
  DFF_X1 OUT2_reg_8_ ( .D(n2546), .CK(CLK), .Q(OUT2[8]), .QN(n3911) );
  DFF_X1 OUT2_reg_6_ ( .D(n2544), .CK(CLK), .Q(OUT2[6]), .QN(n3909) );
  DFF_X1 OUT2_reg_4_ ( .D(n2542), .CK(CLK), .Q(OUT2[4]), .QN(n3907) );
  DFF_X1 OUT2_reg_22_ ( .D(n2560), .CK(CLK), .Q(OUT2[22]), .QN(n3925) );
  DFF_X1 OUT2_reg_20_ ( .D(n2558), .CK(CLK), .Q(OUT2[20]), .QN(n3923) );
  DFF_X1 OUT2_reg_18_ ( .D(n2556), .CK(CLK), .Q(OUT2[18]), .QN(n3921) );
  DFF_X1 OUT2_reg_16_ ( .D(n2554), .CK(CLK), .Q(OUT2[16]), .QN(n3919) );
  DFF_X1 OUT2_reg_14_ ( .D(n2552), .CK(CLK), .Q(OUT2[14]), .QN(n3917) );
  DFF_X1 OUT2_reg_12_ ( .D(n2550), .CK(CLK), .Q(OUT2[12]), .QN(n3915) );
  DFF_X1 OUT1_reg_0_ ( .D(n2506), .CK(CLK), .Q(OUT1[0]), .QN(n3871) );
  DFF_X1 OUT1_reg_31_ ( .D(n2537), .CK(CLK), .Q(OUT1[31]), .QN(n3902) );
  DFF_X1 OUT1_reg_30_ ( .D(n2536), .CK(CLK), .Q(OUT1[30]), .QN(n3901) );
  DFF_X1 OUT1_reg_29_ ( .D(n2535), .CK(CLK), .Q(OUT1[29]), .QN(n3900) );
  DFF_X1 OUT1_reg_28_ ( .D(n2534), .CK(CLK), .Q(OUT1[28]), .QN(n3899) );
  DFF_X1 OUT1_reg_27_ ( .D(n2533), .CK(CLK), .Q(OUT1[27]), .QN(n3898) );
  DFF_X1 OUT1_reg_26_ ( .D(n2532), .CK(CLK), .Q(OUT1[26]), .QN(n3897) );
  DFF_X1 OUT1_reg_25_ ( .D(n2531), .CK(CLK), .Q(OUT1[25]), .QN(n3896) );
  DFF_X1 OUT1_reg_24_ ( .D(n2530), .CK(CLK), .Q(OUT1[24]), .QN(n3895) );
  DFF_X1 OUT1_reg_6_ ( .D(n2512), .CK(CLK), .Q(OUT1[6]), .QN(n3877) );
  DFF_X1 OUT1_reg_5_ ( .D(n2511), .CK(CLK), .Q(OUT1[5]), .QN(n3876) );
  DFF_X1 OUT2_reg_0_ ( .D(n2538), .CK(CLK), .Q(OUT2[0]), .QN(n3903) );
  DFF_X1 OUT2_reg_1_ ( .D(n2539), .CK(CLK), .Q(OUT2[1]), .QN(n3904) );
  DFF_X1 OUT2_reg_2_ ( .D(n2540), .CK(CLK), .Q(OUT2[2]), .QN(n3905) );
  DFF_X1 OUT1_reg_23_ ( .D(n2529), .CK(CLK), .Q(OUT1[23]), .QN(n3894) );
  DFF_X1 OUT1_reg_22_ ( .D(n2528), .CK(CLK), .Q(OUT1[22]), .QN(n3893) );
  DFF_X1 OUT1_reg_21_ ( .D(n2527), .CK(CLK), .Q(OUT1[21]), .QN(n3892) );
  DFF_X1 OUT1_reg_20_ ( .D(n2526), .CK(CLK), .Q(OUT1[20]), .QN(n3891) );
  DFF_X1 OUT1_reg_19_ ( .D(n2525), .CK(CLK), .Q(OUT1[19]), .QN(n3890) );
  DFF_X1 OUT1_reg_18_ ( .D(n2524), .CK(CLK), .Q(OUT1[18]), .QN(n3889) );
  DFF_X1 OUT1_reg_11_ ( .D(n2517), .CK(CLK), .Q(OUT1[11]), .QN(n3882) );
  DFF_X1 OUT1_reg_10_ ( .D(n2516), .CK(CLK), .Q(OUT1[10]), .QN(n3881) );
  DFF_X1 OUT1_reg_7_ ( .D(n2513), .CK(CLK), .Q(OUT1[7]), .QN(n3878) );
  DFF_X1 OUT2_reg_19_ ( .D(n2557), .CK(CLK), .Q(OUT2[19]), .QN(n3922) );
  DFF_X1 OUT2_reg_17_ ( .D(n2555), .CK(CLK), .Q(OUT2[17]), .QN(n3920) );
  DFF_X1 OUT2_reg_15_ ( .D(n2553), .CK(CLK), .Q(OUT2[15]), .QN(n3918) );
  DFF_X1 OUT2_reg_23_ ( .D(n2561), .CK(CLK), .Q(OUT2[23]), .QN(n3926) );
  DFF_X1 OUT2_reg_21_ ( .D(n2559), .CK(CLK), .Q(OUT2[21]), .QN(n3924) );
  DFF_X1 OUT2_reg_13_ ( .D(n2551), .CK(CLK), .Q(OUT2[13]), .QN(n3916) );
  DFF_X1 OUT2_reg_9_ ( .D(n2547), .CK(CLK), .Q(OUT2[9]), .QN(n3912) );
  DFF_X1 OUT2_reg_7_ ( .D(n2545), .CK(CLK), .Q(OUT2[7]), .QN(n3910) );
  DFF_X1 OUT2_reg_5_ ( .D(n2543), .CK(CLK), .Q(OUT2[5]), .QN(n3908) );
  DFF_X1 OUT2_reg_31_ ( .D(n2569), .CK(CLK), .Q(OUT2[31]), .QN(n3934) );
  DFF_X1 OUT2_reg_30_ ( .D(n2568), .CK(CLK), .Q(OUT2[30]), .QN(n3933) );
  DFF_X1 OUT2_reg_29_ ( .D(n2567), .CK(CLK), .Q(OUT2[29]), .QN(n3932) );
  DFF_X1 OUT2_reg_28_ ( .D(n2566), .CK(CLK), .Q(OUT2[28]), .QN(n3931) );
  DFF_X1 OUT2_reg_27_ ( .D(n2565), .CK(CLK), .Q(OUT2[27]), .QN(n3930) );
  DFF_X1 OUT2_reg_26_ ( .D(n2564), .CK(CLK), .Q(OUT2[26]), .QN(n3929) );
  DFF_X1 OUT2_reg_25_ ( .D(n2563), .CK(CLK), .Q(OUT2[25]), .QN(n3928) );
  DFF_X1 OUT2_reg_24_ ( .D(n2562), .CK(CLK), .Q(OUT2[24]), .QN(n3927) );
  DFF_X1 OUT2_reg_11_ ( .D(n2549), .CK(CLK), .Q(OUT2[11]), .QN(n3914) );
  DFF_X2 OUT2_reg_3_ ( .D(n2541), .CK(CLK), .Q(OUT2[3]), .QN(n3906) );
  CLKBUF_X1 U2 ( .A(ADD_RS2[0]), .Z(n1) );
  NOR3_X1 U3 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[3]), .A3(n56), .ZN(n2) );
  CLKBUF_X1 U4 ( .A(n3858), .Z(n3) );
  BUF_X2 U5 ( .A(n1354), .Z(n323) );
  BUF_X2 U6 ( .A(n1353), .Z(n320) );
  BUF_X2 U7 ( .A(n1347), .Z(n309) );
  BUF_X2 U8 ( .A(n1354), .Z(n322) );
  BUF_X2 U9 ( .A(n1353), .Z(n319) );
  BUF_X2 U10 ( .A(n1350), .Z(n315) );
  BUF_X2 U11 ( .A(n1352), .Z(n318) );
  BUF_X2 U12 ( .A(n1343), .Z(n302) );
  BUF_X2 U13 ( .A(n1343), .Z(n301) );
  OAI211_X1 U14 ( .C1(n535), .C2(n305), .A(n1817), .B(n1818), .ZN(n1810) );
  OAI211_X1 U15 ( .C1(n547), .C2(n304), .A(n2117), .B(n2118), .ZN(n2110) );
  BUF_X1 U16 ( .A(n2195), .Z(n457) );
  CLKBUF_X1 U17 ( .A(ADD_RS2[1]), .Z(n4) );
  BUF_X2 U18 ( .A(n1367), .Z(n342) );
  BUF_X2 U19 ( .A(n1367), .Z(n33) );
  BUF_X2 U20 ( .A(n1367), .Z(n34) );
  BUF_X2 U21 ( .A(n1367), .Z(n341) );
  BUF_X2 U22 ( .A(n1367), .Z(n340) );
  CLKBUF_X3 U23 ( .A(n1382), .Z(n5) );
  BUF_X2 U24 ( .A(n1369), .Z(n346) );
  BUF_X2 U25 ( .A(n1369), .Z(n347) );
  CLKBUF_X3 U26 ( .A(n1375), .Z(n356) );
  OR2_X1 U27 ( .A1(n1812), .A2(n1811), .ZN(n6) );
  OR2_X1 U28 ( .A1(n2470), .A2(n2471), .ZN(n7) );
  OR2_X1 U29 ( .A1(n2489), .A2(n2488), .ZN(n8) );
  OR2_X1 U30 ( .A1(n3725), .A2(n3724), .ZN(n9) );
  OR2_X1 U31 ( .A1(n3563), .A2(n3562), .ZN(n10) );
  OR2_X1 U32 ( .A1(n3743), .A2(n3742), .ZN(n11) );
  OR2_X1 U33 ( .A1(n3581), .A2(n3580), .ZN(n12) );
  OR2_X1 U34 ( .A1(n2061), .A2(n2062), .ZN(n13) );
  OR2_X1 U35 ( .A1(n3599), .A2(n3598), .ZN(n14) );
  OR2_X1 U36 ( .A1(n2111), .A2(n2112), .ZN(n15) );
  OR2_X1 U37 ( .A1(n3617), .A2(n3616), .ZN(n16) );
  OR2_X1 U38 ( .A1(n2137), .A2(n2138), .ZN(n17) );
  CLKBUF_X1 U39 ( .A(n2162), .Z(n19) );
  CLKBUF_X3 U40 ( .A(n1350), .Z(n313) );
  BUF_X2 U41 ( .A(n1347), .Z(n307) );
  CLKBUF_X3 U42 ( .A(n1350), .Z(n314) );
  BUF_X2 U43 ( .A(n2206), .Z(n477) );
  CLKBUF_X3 U44 ( .A(n2206), .Z(n476) );
  CLKBUF_X3 U45 ( .A(n2206), .Z(n478) );
  CLKBUF_X1 U46 ( .A(n2143), .Z(n18) );
  BUF_X2 U47 ( .A(n1370), .Z(n349) );
  AND2_X2 U48 ( .A1(ADD_RS2[1]), .A2(n2173), .ZN(n2142) );
  BUF_X1 U49 ( .A(ADD_RS2[3]), .Z(n80) );
  CLKBUF_X3 U50 ( .A(n1363), .Z(n20) );
  CLKBUF_X3 U51 ( .A(n1363), .Z(n21) );
  CLKBUF_X3 U52 ( .A(n1382), .Z(n22) );
  CLKBUF_X3 U53 ( .A(n1382), .Z(n23) );
  CLKBUF_X3 U54 ( .A(n2222), .Z(n24) );
  CLKBUF_X3 U55 ( .A(n2222), .Z(n25) );
  CLKBUF_X1 U56 ( .A(n2149), .Z(n78) );
  CLKBUF_X1 U57 ( .A(n2156), .Z(n26) );
  NOR3_X1 U58 ( .A1(n2469), .A2(n2468), .A3(n7), .ZN(n2467) );
  BUF_X1 U59 ( .A(n2205), .Z(n27) );
  BUF_X1 U60 ( .A(n2205), .Z(n28) );
  BUF_X1 U61 ( .A(n1337), .Z(n29) );
  BUF_X1 U62 ( .A(n1337), .Z(n30) );
  NOR3_X1 U63 ( .A1(n2487), .A2(n2486), .A3(n8), .ZN(n2485) );
  NOR3_X1 U64 ( .A1(n3723), .A2(n3722), .A3(n9), .ZN(n3721) );
  NOR3_X1 U65 ( .A1(n2505), .A2(n2504), .A3(n10), .ZN(n2503) );
  NOR3_X1 U66 ( .A1(n3741), .A2(n3740), .A3(n11), .ZN(n3739) );
  NOR3_X1 U67 ( .A1(n3579), .A2(n3578), .A3(n12), .ZN(n3577) );
  BUF_X1 U68 ( .A(n1362), .Z(n31) );
  BUF_X1 U69 ( .A(n1362), .Z(n32) );
  NOR3_X1 U70 ( .A1(n1809), .A2(n1810), .A3(n6), .ZN(n1808) );
  CLKBUF_X3 U71 ( .A(n1368), .Z(n344) );
  CLKBUF_X2 U72 ( .A(n1368), .Z(n345) );
  CLKBUF_X3 U73 ( .A(n1368), .Z(n343) );
  NOR3_X1 U74 ( .A1(n2059), .A2(n2060), .A3(n13), .ZN(n2058) );
  CLKBUF_X3 U75 ( .A(n1380), .Z(n428) );
  NOR3_X1 U76 ( .A1(n3596), .A2(n3597), .A3(n14), .ZN(n3595) );
  CLKBUF_X3 U77 ( .A(n2216), .Z(n492) );
  NOR3_X1 U78 ( .A1(n2109), .A2(n2110), .A3(n15), .ZN(n2108) );
  NOR3_X1 U79 ( .A1(n3614), .A2(n3615), .A3(n16), .ZN(n3613) );
  CLKBUF_X3 U80 ( .A(n2217), .Z(n496) );
  CLKBUF_X3 U81 ( .A(n2217), .Z(n495) );
  NOR3_X1 U82 ( .A1(n2135), .A2(n2136), .A3(n17), .ZN(n2133) );
  CLKBUF_X3 U83 ( .A(n1380), .Z(n429) );
  BUF_X1 U84 ( .A(n2163), .Z(n35) );
  CLKBUF_X1 U85 ( .A(n3854), .Z(n36) );
  BUF_X2 U86 ( .A(n1377), .Z(n425) );
  BUF_X2 U87 ( .A(n1339), .Z(n228) );
  BUF_X1 U88 ( .A(n1339), .Z(n293) );
  BUF_X1 U89 ( .A(n1377), .Z(n427) );
  BUF_X1 U90 ( .A(n716), .Z(n715) );
  BUF_X1 U91 ( .A(n1347), .Z(n308) );
  BUF_X2 U92 ( .A(n1336), .Z(n222) );
  BUF_X2 U93 ( .A(n1336), .Z(n223) );
  BUF_X2 U94 ( .A(n1360), .Z(n329) );
  BUF_X2 U95 ( .A(n1348), .Z(n310) );
  BUF_X2 U96 ( .A(n1348), .Z(n311) );
  BUF_X2 U97 ( .A(n1365), .Z(n337) );
  BUF_X2 U98 ( .A(n1365), .Z(n338) );
  BUF_X2 U99 ( .A(n1352), .Z(n316) );
  BUF_X2 U100 ( .A(n1375), .Z(n355) );
  BUF_X2 U101 ( .A(n1352), .Z(n317) );
  BUF_X2 U102 ( .A(n1332), .Z(n216) );
  BUF_X2 U103 ( .A(n1332), .Z(n217) );
  BUF_X2 U104 ( .A(n1373), .Z(n352) );
  BUF_X2 U105 ( .A(n1373), .Z(n353) );
  BUF_X2 U106 ( .A(n1334), .Z(n219) );
  BUF_X2 U107 ( .A(n1340), .Z(n295) );
  BUF_X2 U108 ( .A(n1334), .Z(n220) );
  BUF_X2 U109 ( .A(n1340), .Z(n296) );
  BUF_X2 U110 ( .A(n1337), .Z(n225) );
  BUF_X1 U111 ( .A(n1337), .Z(n226) );
  BUF_X2 U112 ( .A(n1359), .Z(n326) );
  BUF_X2 U113 ( .A(n1364), .Z(n334) );
  BUF_X2 U114 ( .A(n1364), .Z(n335) );
  BUF_X2 U115 ( .A(n1344), .Z(n304) );
  BUF_X2 U116 ( .A(n1344), .Z(n305) );
  BUF_X1 U117 ( .A(n1362), .Z(n333) );
  BUF_X1 U118 ( .A(n1362), .Z(n332) );
  BUF_X2 U119 ( .A(n1376), .Z(n422) );
  BUF_X2 U120 ( .A(n1376), .Z(n423) );
  BUF_X1 U121 ( .A(n1362), .Z(n331) );
  BUF_X2 U122 ( .A(n1353), .Z(n321) );
  BUF_X2 U123 ( .A(n1342), .Z(n300) );
  BUF_X1 U124 ( .A(n1336), .Z(n224) );
  BUF_X2 U125 ( .A(n1360), .Z(n330) );
  BUF_X2 U126 ( .A(n1348), .Z(n312) );
  BUF_X2 U127 ( .A(n1365), .Z(n339) );
  BUF_X2 U128 ( .A(n1375), .Z(n421) );
  BUF_X1 U129 ( .A(n1332), .Z(n218) );
  BUF_X2 U130 ( .A(n1373), .Z(n354) );
  BUF_X1 U131 ( .A(n1340), .Z(n297) );
  BUF_X1 U132 ( .A(n1334), .Z(n221) );
  BUF_X2 U133 ( .A(n1380), .Z(n430) );
  BUF_X2 U134 ( .A(n1354), .Z(n324) );
  BUF_X1 U135 ( .A(n1343), .Z(n303) );
  BUF_X1 U136 ( .A(n1337), .Z(n227) );
  BUF_X1 U137 ( .A(n1359), .Z(n327) );
  BUF_X1 U138 ( .A(n1364), .Z(n336) );
  BUF_X1 U139 ( .A(n1369), .Z(n348) );
  BUF_X1 U140 ( .A(n1344), .Z(n306) );
  BUF_X1 U141 ( .A(n594), .Z(n716) );
  BUF_X1 U142 ( .A(n595), .Z(n720) );
  BUF_X1 U143 ( .A(n595), .Z(n721) );
  BUF_X1 U144 ( .A(n595), .Z(n719) );
  BUF_X1 U145 ( .A(n594), .Z(n718) );
  BUF_X1 U146 ( .A(n594), .Z(n717) );
  BUF_X1 U147 ( .A(n597), .Z(n727) );
  BUF_X1 U148 ( .A(n596), .Z(n723) );
  BUF_X1 U149 ( .A(n597), .Z(n726) );
  BUF_X1 U150 ( .A(n597), .Z(n725) );
  BUF_X1 U151 ( .A(n596), .Z(n724) );
  BUF_X1 U152 ( .A(n596), .Z(n722) );
  BUF_X1 U153 ( .A(n598), .Z(n728) );
  BUF_X1 U154 ( .A(n598), .Z(n729) );
  BUF_X2 U155 ( .A(n2192), .Z(n446) );
  BUF_X2 U156 ( .A(n2192), .Z(n447) );
  BUF_X2 U157 ( .A(n2207), .Z(n479) );
  BUF_X2 U158 ( .A(n2197), .Z(n458) );
  BUF_X2 U159 ( .A(n2207), .Z(n480) );
  BUF_X2 U160 ( .A(n2197), .Z(n459) );
  BUF_X2 U161 ( .A(n2203), .Z(n471) );
  BUF_X2 U162 ( .A(n2224), .Z(n510) );
  BUF_X2 U163 ( .A(n2229), .Z(n554) );
  BUF_X2 U164 ( .A(n2214), .Z(n488) );
  BUF_X2 U165 ( .A(n2214), .Z(n489) );
  BUF_X2 U166 ( .A(n2219), .Z(n500) );
  BUF_X2 U167 ( .A(n2219), .Z(n501) );
  BUF_X2 U168 ( .A(n2217), .Z(n494) );
  BUF_X2 U169 ( .A(n2232), .Z(n559) );
  BUF_X2 U170 ( .A(n2232), .Z(n560) );
  BUF_X2 U171 ( .A(n2189), .Z(n440) );
  BUF_X2 U172 ( .A(n2189), .Z(n441) );
  BUF_X2 U173 ( .A(n2194), .Z(n452) );
  BUF_X2 U174 ( .A(n2194), .Z(n453) );
  BUF_X2 U175 ( .A(n2231), .Z(n556) );
  BUF_X2 U176 ( .A(n2231), .Z(n557) );
  BUF_X2 U177 ( .A(n2221), .Z(n503) );
  BUF_X2 U178 ( .A(n2216), .Z(n491) );
  BUF_X2 U179 ( .A(n2226), .Z(n512) );
  BUF_X2 U180 ( .A(n2221), .Z(n504) );
  BUF_X2 U181 ( .A(n2226), .Z(n513) );
  BUF_X1 U182 ( .A(n2205), .Z(n473) );
  BUF_X1 U183 ( .A(n2205), .Z(n474) );
  BUF_X2 U184 ( .A(n2190), .Z(n443) );
  BUF_X2 U185 ( .A(n2195), .Z(n455) );
  BUF_X2 U186 ( .A(n2190), .Z(n444) );
  BUF_X2 U187 ( .A(n2195), .Z(n456) );
  BUF_X2 U188 ( .A(n2208), .Z(n482) );
  BUF_X2 U189 ( .A(n2198), .Z(n461) );
  BUF_X2 U190 ( .A(n2208), .Z(n483) );
  BUF_X2 U191 ( .A(n2193), .Z(n450) );
  BUF_X2 U192 ( .A(n2198), .Z(n462) );
  BUF_X1 U193 ( .A(n2193), .Z(n449) );
  BUF_X2 U194 ( .A(n2202), .Z(n468) );
  BUF_X2 U195 ( .A(n2228), .Z(n551) );
  BUF_X2 U196 ( .A(n2223), .Z(n507) );
  BUF_X2 U197 ( .A(n2218), .Z(n497) );
  BUF_X2 U198 ( .A(n2213), .Z(n485) );
  BUF_X2 U199 ( .A(n2213), .Z(n486) );
  BUF_X2 U200 ( .A(n2218), .Z(n498) );
  BUF_X2 U201 ( .A(n2199), .Z(n464) );
  BUF_X2 U202 ( .A(n2199), .Z(n465) );
  BUF_X2 U203 ( .A(n2227), .Z(n516) );
  BUF_X2 U204 ( .A(n2227), .Z(n549) );
  BUF_X1 U205 ( .A(n2192), .Z(n448) );
  BUF_X1 U206 ( .A(n2197), .Z(n460) );
  BUF_X1 U207 ( .A(n2207), .Z(n481) );
  BUF_X1 U208 ( .A(n2203), .Z(n472) );
  BUF_X1 U209 ( .A(n2224), .Z(n511) );
  BUF_X1 U210 ( .A(n2229), .Z(n555) );
  BUF_X1 U211 ( .A(n2214), .Z(n490) );
  BUF_X1 U212 ( .A(n2219), .Z(n502) );
  BUF_X1 U213 ( .A(n2189), .Z(n442) );
  BUF_X2 U214 ( .A(n2194), .Z(n454) );
  BUF_X2 U215 ( .A(n2231), .Z(n558) );
  BUF_X2 U216 ( .A(n2226), .Z(n514) );
  BUF_X2 U217 ( .A(n2221), .Z(n505) );
  BUF_X2 U218 ( .A(n2216), .Z(n493) );
  BUF_X2 U219 ( .A(n2205), .Z(n475) );
  BUF_X2 U220 ( .A(n2190), .Z(n445) );
  BUF_X1 U221 ( .A(n2202), .Z(n469) );
  BUF_X1 U222 ( .A(n2228), .Z(n552) );
  BUF_X1 U223 ( .A(n2193), .Z(n451) );
  BUF_X1 U224 ( .A(n2208), .Z(n484) );
  BUF_X1 U225 ( .A(n2198), .Z(n463) );
  BUF_X1 U226 ( .A(n2223), .Z(n508) );
  BUF_X1 U227 ( .A(n2218), .Z(n499) );
  BUF_X1 U228 ( .A(n2213), .Z(n487) );
  BUF_X1 U229 ( .A(n2199), .Z(n466) );
  BUF_X1 U230 ( .A(n599), .Z(n597) );
  BUF_X1 U231 ( .A(n599), .Z(n596) );
  BUF_X1 U232 ( .A(n600), .Z(n595) );
  BUF_X1 U233 ( .A(n600), .Z(n594) );
  BUF_X1 U234 ( .A(n599), .Z(n598) );
  BUF_X1 U235 ( .A(n1257), .Z(n201) );
  BUF_X1 U236 ( .A(n1257), .Z(n202) );
  BUF_X1 U237 ( .A(n1222), .Z(n192) );
  BUF_X1 U238 ( .A(n1222), .Z(n193) );
  BUF_X1 U239 ( .A(n1116), .Z(n171) );
  BUF_X1 U240 ( .A(n1116), .Z(n172) );
  BUF_X1 U241 ( .A(n1081), .Z(n162) );
  BUF_X1 U242 ( .A(n1081), .Z(n163) );
  BUF_X1 U243 ( .A(n1012), .Z(n150) );
  BUF_X1 U244 ( .A(n1012), .Z(n151) );
  BUF_X1 U245 ( .A(n979), .Z(n147) );
  BUF_X1 U246 ( .A(n979), .Z(n148) );
  BUF_X1 U247 ( .A(n912), .Z(n138) );
  BUF_X1 U248 ( .A(n912), .Z(n139) );
  BUF_X1 U249 ( .A(n877), .Z(n135) );
  BUF_X1 U250 ( .A(n877), .Z(n136) );
  BUF_X1 U251 ( .A(n1290), .Z(n204) );
  BUF_X1 U252 ( .A(n1290), .Z(n205) );
  BUF_X1 U253 ( .A(n1255), .Z(n198) );
  BUF_X1 U254 ( .A(n1255), .Z(n199) );
  BUF_X1 U255 ( .A(n1254), .Z(n195) );
  BUF_X1 U256 ( .A(n1254), .Z(n196) );
  BUF_X1 U257 ( .A(n1188), .Z(n189) );
  BUF_X1 U258 ( .A(n1188), .Z(n190) );
  BUF_X1 U259 ( .A(n1185), .Z(n186) );
  BUF_X1 U260 ( .A(n1185), .Z(n187) );
  BUF_X1 U261 ( .A(n1183), .Z(n183) );
  BUF_X1 U262 ( .A(n1183), .Z(n184) );
  BUF_X1 U263 ( .A(n1182), .Z(n180) );
  BUF_X1 U264 ( .A(n1182), .Z(n181) );
  BUF_X1 U265 ( .A(n1181), .Z(n177) );
  BUF_X1 U266 ( .A(n1181), .Z(n178) );
  BUF_X1 U267 ( .A(n1149), .Z(n174) );
  BUF_X1 U268 ( .A(n1149), .Z(n175) );
  BUF_X1 U269 ( .A(n1114), .Z(n168) );
  BUF_X1 U270 ( .A(n1114), .Z(n169) );
  BUF_X1 U271 ( .A(n1113), .Z(n165) );
  BUF_X1 U272 ( .A(n1113), .Z(n166) );
  BUF_X1 U273 ( .A(n1047), .Z(n159) );
  BUF_X1 U274 ( .A(n1047), .Z(n160) );
  BUF_X1 U275 ( .A(n1045), .Z(n156) );
  BUF_X1 U276 ( .A(n1045), .Z(n157) );
  BUF_X1 U277 ( .A(n1044), .Z(n153) );
  BUF_X1 U278 ( .A(n1044), .Z(n154) );
  BUF_X1 U279 ( .A(n977), .Z(n144) );
  BUF_X1 U280 ( .A(n977), .Z(n145) );
  BUF_X1 U281 ( .A(n976), .Z(n141) );
  BUF_X1 U282 ( .A(n976), .Z(n142) );
  BUF_X1 U283 ( .A(n871), .Z(n132) );
  BUF_X1 U284 ( .A(n871), .Z(n133) );
  BUF_X1 U285 ( .A(n869), .Z(n129) );
  BUF_X1 U286 ( .A(n869), .Z(n130) );
  BUF_X1 U287 ( .A(n804), .Z(n126) );
  BUF_X1 U288 ( .A(n804), .Z(n127) );
  BUF_X1 U289 ( .A(n770), .Z(n123) );
  BUF_X1 U290 ( .A(n770), .Z(n124) );
  BUF_X1 U291 ( .A(n767), .Z(n120) );
  BUF_X1 U292 ( .A(n767), .Z(n121) );
  BUF_X1 U293 ( .A(n765), .Z(n117) );
  BUF_X1 U294 ( .A(n765), .Z(n118) );
  BUF_X1 U295 ( .A(n731), .Z(n114) );
  BUF_X1 U296 ( .A(n731), .Z(n115) );
  BUF_X2 U297 ( .A(n2183), .Z(n434) );
  BUF_X2 U298 ( .A(n2183), .Z(n435) );
  BUF_X2 U299 ( .A(n1324), .Z(n207) );
  BUF_X2 U300 ( .A(n1324), .Z(n208) );
  BUF_X2 U301 ( .A(n2181), .Z(n431) );
  BUF_X2 U302 ( .A(n2181), .Z(n432) );
  BUF_X1 U303 ( .A(n1257), .Z(n203) );
  BUF_X1 U304 ( .A(n1222), .Z(n194) );
  BUF_X1 U305 ( .A(n1116), .Z(n173) );
  BUF_X1 U306 ( .A(n1081), .Z(n164) );
  BUF_X1 U307 ( .A(n1012), .Z(n152) );
  BUF_X1 U308 ( .A(n979), .Z(n149) );
  BUF_X1 U309 ( .A(n912), .Z(n140) );
  BUF_X1 U310 ( .A(n877), .Z(n137) );
  BUF_X1 U311 ( .A(n1290), .Z(n206) );
  BUF_X1 U312 ( .A(n1255), .Z(n200) );
  BUF_X1 U313 ( .A(n1254), .Z(n197) );
  BUF_X1 U314 ( .A(n1188), .Z(n191) );
  BUF_X1 U315 ( .A(n1185), .Z(n188) );
  BUF_X1 U316 ( .A(n1183), .Z(n185) );
  BUF_X1 U317 ( .A(n1182), .Z(n182) );
  BUF_X1 U318 ( .A(n1181), .Z(n179) );
  BUF_X1 U319 ( .A(n1149), .Z(n176) );
  BUF_X1 U320 ( .A(n1114), .Z(n170) );
  BUF_X1 U321 ( .A(n1113), .Z(n167) );
  BUF_X1 U322 ( .A(n1047), .Z(n161) );
  BUF_X1 U323 ( .A(n767), .Z(n122) );
  BUF_X1 U324 ( .A(n765), .Z(n119) );
  BUF_X1 U325 ( .A(n731), .Z(n116) );
  BUF_X1 U326 ( .A(n1045), .Z(n158) );
  BUF_X1 U327 ( .A(n1044), .Z(n155) );
  BUF_X1 U328 ( .A(n977), .Z(n146) );
  BUF_X1 U329 ( .A(n976), .Z(n143) );
  BUF_X1 U330 ( .A(n871), .Z(n134) );
  BUF_X1 U331 ( .A(n869), .Z(n131) );
  BUF_X1 U332 ( .A(n804), .Z(n128) );
  BUF_X1 U333 ( .A(n770), .Z(n125) );
  BUF_X1 U334 ( .A(n2183), .Z(n436) );
  BUF_X1 U335 ( .A(n1326), .Z(n212) );
  BUF_X1 U336 ( .A(n2181), .Z(n433) );
  BUF_X1 U337 ( .A(n1324), .Z(n209) );
  BUF_X1 U338 ( .A(RST), .Z(n599) );
  BUF_X1 U339 ( .A(RST), .Z(n600) );
  BUF_X1 U340 ( .A(n2184), .Z(n437) );
  BUF_X1 U341 ( .A(n1327), .Z(n213) );
  BUF_X1 U342 ( .A(n2184), .Z(n438) );
  BUF_X1 U343 ( .A(n1327), .Z(n214) );
  BUF_X1 U344 ( .A(n2184), .Z(n439) );
  BUF_X1 U345 ( .A(n1327), .Z(n215) );
  INV_X1 U346 ( .A(DATAIN[2]), .ZN(n564) );
  INV_X1 U347 ( .A(DATAIN[4]), .ZN(n566) );
  INV_X1 U348 ( .A(DATAIN[5]), .ZN(n567) );
  INV_X1 U349 ( .A(DATAIN[6]), .ZN(n568) );
  INV_X1 U350 ( .A(DATAIN[7]), .ZN(n569) );
  INV_X1 U351 ( .A(DATAIN[8]), .ZN(n570) );
  INV_X1 U352 ( .A(DATAIN[10]), .ZN(n572) );
  INV_X1 U353 ( .A(DATAIN[11]), .ZN(n573) );
  INV_X1 U354 ( .A(DATAIN[12]), .ZN(n574) );
  INV_X1 U355 ( .A(DATAIN[13]), .ZN(n575) );
  INV_X1 U356 ( .A(DATAIN[14]), .ZN(n576) );
  INV_X1 U357 ( .A(DATAIN[15]), .ZN(n577) );
  INV_X1 U358 ( .A(DATAIN[16]), .ZN(n578) );
  INV_X1 U359 ( .A(DATAIN[17]), .ZN(n579) );
  INV_X1 U360 ( .A(DATAIN[18]), .ZN(n580) );
  INV_X1 U361 ( .A(DATAIN[19]), .ZN(n581) );
  INV_X1 U362 ( .A(DATAIN[20]), .ZN(n582) );
  INV_X1 U363 ( .A(DATAIN[21]), .ZN(n583) );
  INV_X1 U364 ( .A(DATAIN[22]), .ZN(n584) );
  INV_X1 U365 ( .A(DATAIN[23]), .ZN(n585) );
  INV_X1 U366 ( .A(DATAIN[24]), .ZN(n586) );
  INV_X1 U367 ( .A(DATAIN[25]), .ZN(n587) );
  INV_X1 U368 ( .A(DATAIN[26]), .ZN(n588) );
  INV_X1 U369 ( .A(DATAIN[27]), .ZN(n589) );
  INV_X1 U370 ( .A(DATAIN[28]), .ZN(n590) );
  INV_X1 U371 ( .A(DATAIN[29]), .ZN(n591) );
  INV_X1 U372 ( .A(DATAIN[30]), .ZN(n592) );
  INV_X1 U373 ( .A(DATAIN[31]), .ZN(n593) );
  INV_X1 U374 ( .A(DATAIN[0]), .ZN(n562) );
  INV_X1 U375 ( .A(DATAIN[1]), .ZN(n563) );
  INV_X1 U376 ( .A(DATAIN[3]), .ZN(n565) );
  INV_X1 U377 ( .A(DATAIN[9]), .ZN(n571) );
  OR2_X1 U378 ( .A1(n3815), .A2(n3814), .ZN(n37) );
  OR2_X1 U379 ( .A1(n3797), .A2(n3796), .ZN(n38) );
  OR2_X1 U380 ( .A1(n3779), .A2(n3778), .ZN(n39) );
  OR2_X1 U381 ( .A1(n2037), .A2(n2036), .ZN(n40) );
  OR2_X1 U382 ( .A1(n1987), .A2(n1986), .ZN(n41) );
  OR2_X1 U383 ( .A1(n1937), .A2(n1936), .ZN(n42) );
  OR2_X1 U384 ( .A1(n1887), .A2(n1886), .ZN(n43) );
  OR2_X1 U385 ( .A1(n1837), .A2(n1836), .ZN(n44) );
  OR2_X1 U386 ( .A1(n1787), .A2(n1786), .ZN(n45) );
  OR2_X1 U387 ( .A1(n1737), .A2(n1736), .ZN(n46) );
  OR2_X1 U388 ( .A1(n1687), .A2(n1686), .ZN(n47) );
  OR2_X1 U389 ( .A1(n1637), .A2(n1636), .ZN(n48) );
  OR2_X1 U390 ( .A1(n1587), .A2(n1586), .ZN(n49) );
  OR2_X1 U391 ( .A1(n2087), .A2(n2086), .ZN(n50) );
  OR2_X1 U392 ( .A1(n3761), .A2(n3760), .ZN(n51) );
  OR2_X1 U393 ( .A1(n3689), .A2(n3688), .ZN(n52) );
  OR2_X1 U394 ( .A1(n3671), .A2(n3670), .ZN(n53) );
  CLKBUF_X1 U395 ( .A(n2168), .Z(n79) );
  AND3_X1 U396 ( .A1(ADD_RS1[0]), .A2(n56), .A3(ADD_RS1[3]), .ZN(n3855) );
  BUF_X1 U397 ( .A(n2141), .Z(n54) );
  INV_X1 U398 ( .A(ADD_RS1[4]), .ZN(n55) );
  INV_X1 U399 ( .A(ADD_RS1[4]), .ZN(n56) );
  CLKBUF_X1 U400 ( .A(ADD_RS1[2]), .Z(n57) );
  CLKBUF_X1 U401 ( .A(n2), .Z(n58) );
  NAND2_X1 U402 ( .A1(n424), .A2(n739), .ZN(n59) );
  NAND2_X1 U403 ( .A1(n426), .A2(n3958), .ZN(n60) );
  INV_X1 U404 ( .A(n1580), .ZN(n61) );
  AND3_X1 U405 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n1571) );
  NAND2_X1 U406 ( .A1(n424), .A2(n741), .ZN(n62) );
  NAND2_X1 U407 ( .A1(n426), .A2(n3956), .ZN(n63) );
  INV_X1 U408 ( .A(n1630), .ZN(n64) );
  AND3_X1 U409 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n1621) );
  NAND2_X1 U410 ( .A1(n424), .A2(n743), .ZN(n65) );
  NAND2_X1 U411 ( .A1(n426), .A2(n3954), .ZN(n66) );
  INV_X1 U412 ( .A(n1680), .ZN(n67) );
  AND3_X1 U413 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n1671) );
  NAND2_X1 U414 ( .A1(n424), .A2(n745), .ZN(n68) );
  NAND2_X1 U415 ( .A1(n426), .A2(n3952), .ZN(n69) );
  INV_X1 U416 ( .A(n1730), .ZN(n70) );
  AND3_X1 U417 ( .A1(n68), .A2(n69), .A3(n70), .ZN(n1721) );
  NAND2_X1 U418 ( .A1(n424), .A2(n747), .ZN(n71) );
  NAND2_X1 U419 ( .A1(n426), .A2(n3950), .ZN(n72) );
  INV_X1 U420 ( .A(n1780), .ZN(n73) );
  AND3_X1 U421 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n1771) );
  NAND2_X1 U422 ( .A1(n424), .A2(n749), .ZN(n74) );
  NAND2_X1 U423 ( .A1(n426), .A2(n3948), .ZN(n75) );
  INV_X1 U424 ( .A(n1830), .ZN(n76) );
  AND3_X1 U425 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n1821) );
  BUF_X2 U426 ( .A(n1376), .Z(n424) );
  BUF_X2 U427 ( .A(n1377), .Z(n426) );
  CLKBUF_X1 U428 ( .A(n1339), .Z(n294) );
  CLKBUF_X1 U429 ( .A(n2149), .Z(n85) );
  INV_X1 U430 ( .A(ADD_RS2[0]), .ZN(n77) );
  BUF_X1 U431 ( .A(n1370), .Z(n350) );
  BUF_X1 U432 ( .A(n1370), .Z(n351) );
  AND2_X1 U433 ( .A1(n325), .A2(n4194), .ZN(n81) );
  AND2_X1 U434 ( .A1(n328), .A2(n4226), .ZN(n82) );
  NOR3_X1 U435 ( .A1(n81), .A2(n82), .A3(n2075), .ZN(n2074) );
  BUF_X2 U436 ( .A(n1359), .Z(n325) );
  BUF_X2 U437 ( .A(n1360), .Z(n328) );
  INV_X1 U438 ( .A(ADD_RS1[0]), .ZN(n83) );
  INV_X1 U439 ( .A(ADD_RS1[0]), .ZN(n84) );
  CLKBUF_X2 U440 ( .A(n2232), .Z(n561) );
  CLKBUF_X2 U441 ( .A(n2227), .Z(n515) );
  AND2_X1 U442 ( .A1(ADD_RS2[2]), .A2(ADD_RS2[1]), .ZN(n2145) );
  NOR3_X1 U443 ( .A1(n77), .A2(ADD_RS2[4]), .A3(ADD_RS2[3]), .ZN(n2168) );
  INV_X1 U444 ( .A(ADD_RS2[4]), .ZN(n86) );
  NOR3_X1 U445 ( .A1(n1584), .A2(n1585), .A3(n49), .ZN(n1583) );
  NOR3_X1 U446 ( .A1(n1634), .A2(n1635), .A3(n48), .ZN(n1633) );
  NOR3_X1 U447 ( .A1(n1684), .A2(n1685), .A3(n47), .ZN(n1683) );
  NOR3_X1 U448 ( .A1(n1734), .A2(n1735), .A3(n46), .ZN(n1733) );
  NOR3_X1 U449 ( .A1(n1784), .A2(n1785), .A3(n45), .ZN(n1783) );
  NOR3_X1 U450 ( .A1(n1834), .A2(n1835), .A3(n44), .ZN(n1833) );
  NOR3_X1 U451 ( .A1(n1884), .A2(n1885), .A3(n43), .ZN(n1883) );
  NOR3_X1 U452 ( .A1(n1934), .A2(n1935), .A3(n42), .ZN(n1933) );
  NOR3_X1 U453 ( .A1(n1984), .A2(n1985), .A3(n41), .ZN(n1983) );
  NOR3_X1 U454 ( .A1(n2034), .A2(n2035), .A3(n40), .ZN(n2033) );
  AND2_X1 U455 ( .A1(n346), .A2(n799), .ZN(n87) );
  AND2_X1 U456 ( .A1(n349), .A2(n833), .ZN(n88) );
  NOR3_X1 U457 ( .A1(n87), .A2(n88), .A3(n2102), .ZN(n2097) );
  NOR3_X1 U458 ( .A1(n2085), .A2(n2084), .A3(n50), .ZN(n2083) );
  AND2_X1 U459 ( .A1(n346), .A2(n800), .ZN(n89) );
  AND2_X1 U460 ( .A1(n349), .A2(n834), .ZN(n90) );
  NOR3_X1 U461 ( .A1(n89), .A2(n90), .A3(n2127), .ZN(n2122) );
  AND2_X1 U462 ( .A1(n550), .A2(n762), .ZN(n91) );
  AND2_X1 U463 ( .A1(n553), .A2(n3935), .ZN(n92) );
  NOR3_X1 U464 ( .A1(n91), .A2(n92), .A3(n3860), .ZN(n3849) );
  BUF_X2 U465 ( .A(n2228), .Z(n550) );
  BUF_X2 U466 ( .A(n2229), .Z(n553) );
  AND2_X1 U467 ( .A1(n346), .A2(n801), .ZN(n93) );
  AND2_X1 U468 ( .A1(n349), .A2(n835), .ZN(n94) );
  NOR3_X1 U469 ( .A1(n93), .A2(n94), .A3(n2165), .ZN(n2158) );
  AND2_X1 U470 ( .A1(n506), .A2(n790), .ZN(n95) );
  AND2_X1 U471 ( .A1(n509), .A2(n824), .ZN(n96) );
  NOR3_X1 U472 ( .A1(n95), .A2(n96), .A3(n3647), .ZN(n3642) );
  AND2_X1 U473 ( .A1(n506), .A2(n791), .ZN(n97) );
  AND2_X1 U474 ( .A1(n509), .A2(n825), .ZN(n98) );
  NOR3_X1 U475 ( .A1(n97), .A2(n98), .A3(n3665), .ZN(n3660) );
  NOR3_X1 U476 ( .A1(n3668), .A2(n3669), .A3(n53), .ZN(n3667) );
  AND2_X1 U477 ( .A1(n506), .A2(n793), .ZN(n99) );
  AND2_X1 U478 ( .A1(n509), .A2(n827), .ZN(n100) );
  NOR3_X1 U479 ( .A1(n99), .A2(n100), .A3(n3701), .ZN(n3696) );
  NOR3_X1 U480 ( .A1(n3686), .A2(n3687), .A3(n52), .ZN(n3685) );
  AND2_X1 U481 ( .A1(n506), .A2(n794), .ZN(n101) );
  AND2_X1 U482 ( .A1(n509), .A2(n828), .ZN(n102) );
  NOR3_X1 U483 ( .A1(n101), .A2(n102), .A3(n3719), .ZN(n3714) );
  AND2_X1 U484 ( .A1(n506), .A2(n795), .ZN(n103) );
  AND2_X1 U485 ( .A1(n509), .A2(n829), .ZN(n104) );
  NOR3_X1 U486 ( .A1(n103), .A2(n104), .A3(n3737), .ZN(n3732) );
  AND2_X1 U487 ( .A1(n506), .A2(n796), .ZN(n105) );
  AND2_X1 U488 ( .A1(n509), .A2(n830), .ZN(n106) );
  NOR3_X1 U489 ( .A1(n105), .A2(n106), .A3(n3755), .ZN(n3750) );
  NOR3_X1 U490 ( .A1(n3758), .A2(n3759), .A3(n51), .ZN(n3757) );
  AND2_X2 U491 ( .A1(ADD_RS1[2]), .A2(ADD_RS1[1]), .ZN(n3840) );
  NOR3_X1 U492 ( .A1(n3776), .A2(n3777), .A3(n39), .ZN(n3775) );
  AND2_X1 U493 ( .A1(n506), .A2(n799), .ZN(n107) );
  AND2_X1 U494 ( .A1(n509), .A2(n833), .ZN(n108) );
  NOR3_X1 U495 ( .A1(n107), .A2(n108), .A3(n3809), .ZN(n3804) );
  NOR3_X1 U496 ( .A1(n3794), .A2(n3795), .A3(n38), .ZN(n3793) );
  NOR3_X1 U497 ( .A1(n3812), .A2(n3813), .A3(n37), .ZN(n3811) );
  AND2_X1 U498 ( .A1(n506), .A2(n801), .ZN(n109) );
  AND2_X1 U499 ( .A1(n509), .A2(n835), .ZN(n110) );
  NOR3_X1 U500 ( .A1(n109), .A2(n110), .A3(n3857), .ZN(n3850) );
  BUF_X2 U501 ( .A(n2223), .Z(n506) );
  BUF_X2 U502 ( .A(n2224), .Z(n509) );
  AND2_X1 U503 ( .A1(n467), .A2(n1180), .ZN(n111) );
  AND2_X1 U504 ( .A1(n470), .A2(n4127), .ZN(n112) );
  NOR3_X1 U505 ( .A1(n111), .A2(n112), .A3(n3847), .ZN(n3846) );
  NOR2_X1 U506 ( .A1(n3861), .A2(ADD_RS1[1]), .ZN(n113) );
  BUF_X2 U507 ( .A(n2202), .Z(n467) );
  BUF_X2 U508 ( .A(n2203), .Z(n470) );
  CLKBUF_X3 U509 ( .A(n1326), .Z(n210) );
  CLKBUF_X3 U510 ( .A(n1326), .Z(n211) );
  CLKBUF_X3 U511 ( .A(n1342), .Z(n298) );
  CLKBUF_X3 U512 ( .A(n1342), .Z(n299) );
  CLKBUF_X1 U513 ( .A(n729), .Z(n601) );
  CLKBUF_X1 U514 ( .A(n729), .Z(n602) );
  CLKBUF_X1 U515 ( .A(n729), .Z(n603) );
  CLKBUF_X1 U516 ( .A(n729), .Z(n604) );
  CLKBUF_X1 U517 ( .A(n729), .Z(n605) );
  CLKBUF_X1 U518 ( .A(n728), .Z(n606) );
  CLKBUF_X1 U519 ( .A(n728), .Z(n607) );
  CLKBUF_X1 U520 ( .A(n728), .Z(n608) );
  CLKBUF_X1 U521 ( .A(n728), .Z(n609) );
  CLKBUF_X1 U522 ( .A(n728), .Z(n610) );
  CLKBUF_X1 U523 ( .A(n728), .Z(n611) );
  CLKBUF_X1 U524 ( .A(n727), .Z(n612) );
  CLKBUF_X1 U525 ( .A(n727), .Z(n645) );
  CLKBUF_X1 U526 ( .A(n727), .Z(n646) );
  CLKBUF_X1 U527 ( .A(n727), .Z(n647) );
  CLKBUF_X1 U528 ( .A(n727), .Z(n648) );
  CLKBUF_X1 U529 ( .A(n727), .Z(n649) );
  CLKBUF_X1 U530 ( .A(n726), .Z(n650) );
  CLKBUF_X1 U531 ( .A(n726), .Z(n651) );
  CLKBUF_X1 U532 ( .A(n726), .Z(n652) );
  CLKBUF_X1 U533 ( .A(n726), .Z(n653) );
  CLKBUF_X1 U534 ( .A(n726), .Z(n654) );
  CLKBUF_X1 U535 ( .A(n726), .Z(n655) );
  CLKBUF_X1 U536 ( .A(n725), .Z(n656) );
  CLKBUF_X1 U537 ( .A(n725), .Z(n657) );
  CLKBUF_X1 U538 ( .A(n725), .Z(n658) );
  CLKBUF_X1 U539 ( .A(n725), .Z(n659) );
  CLKBUF_X1 U540 ( .A(n725), .Z(n660) );
  CLKBUF_X1 U541 ( .A(n725), .Z(n661) );
  CLKBUF_X1 U542 ( .A(n724), .Z(n662) );
  CLKBUF_X1 U543 ( .A(n724), .Z(n663) );
  CLKBUF_X1 U544 ( .A(n724), .Z(n664) );
  CLKBUF_X1 U545 ( .A(n724), .Z(n665) );
  CLKBUF_X1 U546 ( .A(n724), .Z(n666) );
  CLKBUF_X1 U547 ( .A(n724), .Z(n667) );
  CLKBUF_X1 U548 ( .A(n723), .Z(n668) );
  CLKBUF_X1 U549 ( .A(n723), .Z(n669) );
  CLKBUF_X1 U550 ( .A(n723), .Z(n670) );
  CLKBUF_X1 U551 ( .A(n723), .Z(n671) );
  CLKBUF_X1 U552 ( .A(n723), .Z(n672) );
  CLKBUF_X1 U553 ( .A(n723), .Z(n673) );
  CLKBUF_X1 U554 ( .A(n722), .Z(n674) );
  CLKBUF_X1 U555 ( .A(n722), .Z(n675) );
  CLKBUF_X1 U556 ( .A(n722), .Z(n676) );
  CLKBUF_X1 U557 ( .A(n722), .Z(n677) );
  CLKBUF_X1 U558 ( .A(n722), .Z(n678) );
  CLKBUF_X1 U559 ( .A(n722), .Z(n679) );
  CLKBUF_X1 U560 ( .A(n721), .Z(n680) );
  CLKBUF_X1 U561 ( .A(n721), .Z(n681) );
  CLKBUF_X1 U562 ( .A(n721), .Z(n682) );
  CLKBUF_X1 U563 ( .A(n721), .Z(n683) );
  CLKBUF_X1 U564 ( .A(n721), .Z(n684) );
  CLKBUF_X1 U565 ( .A(n721), .Z(n685) );
  CLKBUF_X1 U566 ( .A(n720), .Z(n686) );
  CLKBUF_X1 U567 ( .A(n720), .Z(n687) );
  CLKBUF_X1 U568 ( .A(n720), .Z(n688) );
  CLKBUF_X1 U569 ( .A(n720), .Z(n689) );
  CLKBUF_X1 U570 ( .A(n720), .Z(n690) );
  CLKBUF_X1 U571 ( .A(n720), .Z(n691) );
  CLKBUF_X1 U572 ( .A(n719), .Z(n692) );
  CLKBUF_X1 U573 ( .A(n719), .Z(n693) );
  CLKBUF_X1 U574 ( .A(n719), .Z(n694) );
  CLKBUF_X1 U575 ( .A(n719), .Z(n695) );
  CLKBUF_X1 U576 ( .A(n719), .Z(n696) );
  CLKBUF_X1 U577 ( .A(n719), .Z(n697) );
  CLKBUF_X1 U578 ( .A(n718), .Z(n698) );
  CLKBUF_X1 U579 ( .A(n718), .Z(n699) );
  CLKBUF_X1 U580 ( .A(n718), .Z(n700) );
  CLKBUF_X1 U581 ( .A(n718), .Z(n701) );
  CLKBUF_X1 U582 ( .A(n718), .Z(n702) );
  CLKBUF_X1 U583 ( .A(n718), .Z(n703) );
  CLKBUF_X1 U584 ( .A(n717), .Z(n704) );
  CLKBUF_X1 U585 ( .A(n717), .Z(n705) );
  CLKBUF_X1 U586 ( .A(n717), .Z(n706) );
  CLKBUF_X1 U587 ( .A(n717), .Z(n707) );
  CLKBUF_X1 U588 ( .A(n717), .Z(n708) );
  CLKBUF_X1 U589 ( .A(n717), .Z(n709) );
  CLKBUF_X1 U590 ( .A(n716), .Z(n710) );
  CLKBUF_X1 U591 ( .A(n716), .Z(n711) );
  CLKBUF_X1 U592 ( .A(n716), .Z(n712) );
  CLKBUF_X1 U593 ( .A(n716), .Z(n713) );
  CLKBUF_X1 U594 ( .A(n716), .Z(n714) );
  MUX2_X1 U595 ( .A(n730), .B(DATAIN[31]), .S(n116), .Z(n3561) );
  MUX2_X1 U596 ( .A(n732), .B(DATAIN[30]), .S(n116), .Z(n3560) );
  MUX2_X1 U597 ( .A(n733), .B(DATAIN[29]), .S(n116), .Z(n3559) );
  MUX2_X1 U598 ( .A(n734), .B(DATAIN[28]), .S(n116), .Z(n3558) );
  MUX2_X1 U599 ( .A(n735), .B(DATAIN[27]), .S(n116), .Z(n3557) );
  MUX2_X1 U600 ( .A(n736), .B(DATAIN[26]), .S(n116), .Z(n3556) );
  MUX2_X1 U601 ( .A(n737), .B(DATAIN[25]), .S(n116), .Z(n3555) );
  MUX2_X1 U602 ( .A(n738), .B(DATAIN[24]), .S(n116), .Z(n3554) );
  MUX2_X1 U603 ( .A(n739), .B(DATAIN[23]), .S(n115), .Z(n3553) );
  MUX2_X1 U604 ( .A(n740), .B(DATAIN[22]), .S(n115), .Z(n3552) );
  MUX2_X1 U605 ( .A(n741), .B(DATAIN[21]), .S(n115), .Z(n3551) );
  MUX2_X1 U606 ( .A(n742), .B(DATAIN[20]), .S(n115), .Z(n3550) );
  MUX2_X1 U607 ( .A(n743), .B(DATAIN[19]), .S(n115), .Z(n3549) );
  MUX2_X1 U608 ( .A(n744), .B(DATAIN[18]), .S(n115), .Z(n3548) );
  MUX2_X1 U609 ( .A(n745), .B(DATAIN[17]), .S(n115), .Z(n3547) );
  MUX2_X1 U610 ( .A(n746), .B(DATAIN[16]), .S(n115), .Z(n3546) );
  MUX2_X1 U611 ( .A(n747), .B(DATAIN[15]), .S(n115), .Z(n3545) );
  MUX2_X1 U612 ( .A(n748), .B(DATAIN[14]), .S(n115), .Z(n3544) );
  MUX2_X1 U613 ( .A(n749), .B(DATAIN[13]), .S(n115), .Z(n3543) );
  MUX2_X1 U614 ( .A(n750), .B(DATAIN[12]), .S(n115), .Z(n3542) );
  MUX2_X1 U615 ( .A(n751), .B(DATAIN[11]), .S(n114), .Z(n3541) );
  MUX2_X1 U616 ( .A(n752), .B(DATAIN[10]), .S(n114), .Z(n3540) );
  MUX2_X1 U617 ( .A(n753), .B(DATAIN[9]), .S(n114), .Z(n3539) );
  MUX2_X1 U618 ( .A(n754), .B(DATAIN[8]), .S(n114), .Z(n3538) );
  MUX2_X1 U619 ( .A(n755), .B(DATAIN[7]), .S(n114), .Z(n3537) );
  MUX2_X1 U620 ( .A(n756), .B(DATAIN[6]), .S(n114), .Z(n3536) );
  MUX2_X1 U621 ( .A(n757), .B(DATAIN[5]), .S(n114), .Z(n3535) );
  MUX2_X1 U622 ( .A(n758), .B(DATAIN[4]), .S(n114), .Z(n3534) );
  MUX2_X1 U623 ( .A(n759), .B(DATAIN[3]), .S(n114), .Z(n3533) );
  MUX2_X1 U624 ( .A(n760), .B(DATAIN[2]), .S(n114), .Z(n3532) );
  MUX2_X1 U625 ( .A(n761), .B(DATAIN[1]), .S(n114), .Z(n3531) );
  MUX2_X1 U626 ( .A(n762), .B(DATAIN[0]), .S(n114), .Z(n3530) );
  AND2_X1 U627 ( .A1(n763), .A2(n764), .ZN(n731) );
  MUX2_X1 U628 ( .A(n4446), .B(DATAIN[31]), .S(n119), .Z(n3529) );
  MUX2_X1 U629 ( .A(n4445), .B(DATAIN[30]), .S(n119), .Z(n3528) );
  MUX2_X1 U630 ( .A(n4444), .B(DATAIN[29]), .S(n119), .Z(n3527) );
  MUX2_X1 U631 ( .A(n4443), .B(DATAIN[28]), .S(n119), .Z(n3526) );
  MUX2_X1 U632 ( .A(n4442), .B(DATAIN[27]), .S(n119), .Z(n3525) );
  MUX2_X1 U633 ( .A(n4441), .B(DATAIN[26]), .S(n119), .Z(n3524) );
  MUX2_X1 U634 ( .A(n4440), .B(DATAIN[25]), .S(n119), .Z(n3523) );
  MUX2_X1 U635 ( .A(n4439), .B(DATAIN[24]), .S(n119), .Z(n3522) );
  MUX2_X1 U636 ( .A(n4438), .B(DATAIN[23]), .S(n118), .Z(n3521) );
  MUX2_X1 U637 ( .A(n4437), .B(DATAIN[22]), .S(n118), .Z(n3520) );
  MUX2_X1 U638 ( .A(n4436), .B(DATAIN[21]), .S(n118), .Z(n3519) );
  MUX2_X1 U639 ( .A(n4435), .B(DATAIN[20]), .S(n118), .Z(n3518) );
  MUX2_X1 U640 ( .A(n4434), .B(DATAIN[19]), .S(n118), .Z(n3517) );
  MUX2_X1 U641 ( .A(n4433), .B(DATAIN[18]), .S(n118), .Z(n3516) );
  MUX2_X1 U642 ( .A(n4432), .B(DATAIN[17]), .S(n118), .Z(n3515) );
  MUX2_X1 U643 ( .A(n4431), .B(DATAIN[16]), .S(n118), .Z(n3514) );
  MUX2_X1 U644 ( .A(n4430), .B(DATAIN[15]), .S(n118), .Z(n3513) );
  MUX2_X1 U645 ( .A(n4429), .B(DATAIN[14]), .S(n118), .Z(n3512) );
  MUX2_X1 U646 ( .A(n4428), .B(DATAIN[13]), .S(n118), .Z(n3511) );
  MUX2_X1 U647 ( .A(n4427), .B(DATAIN[12]), .S(n118), .Z(n3510) );
  MUX2_X1 U648 ( .A(n4426), .B(DATAIN[11]), .S(n117), .Z(n3509) );
  MUX2_X1 U649 ( .A(n4425), .B(DATAIN[10]), .S(n117), .Z(n3508) );
  MUX2_X1 U650 ( .A(n4424), .B(DATAIN[9]), .S(n117), .Z(n3507) );
  MUX2_X1 U651 ( .A(n4423), .B(DATAIN[8]), .S(n117), .Z(n3506) );
  MUX2_X1 U652 ( .A(n4422), .B(DATAIN[7]), .S(n117), .Z(n3505) );
  MUX2_X1 U653 ( .A(n4421), .B(DATAIN[6]), .S(n117), .Z(n3504) );
  MUX2_X1 U654 ( .A(n4420), .B(DATAIN[5]), .S(n117), .Z(n3503) );
  MUX2_X1 U655 ( .A(n4419), .B(DATAIN[4]), .S(n117), .Z(n3502) );
  MUX2_X1 U656 ( .A(n4418), .B(DATAIN[3]), .S(n117), .Z(n3501) );
  MUX2_X1 U657 ( .A(n4417), .B(DATAIN[2]), .S(n117), .Z(n3500) );
  MUX2_X1 U658 ( .A(n4416), .B(DATAIN[1]), .S(n117), .Z(n3499) );
  MUX2_X1 U659 ( .A(n4415), .B(DATAIN[0]), .S(n117), .Z(n3498) );
  AND2_X1 U660 ( .A1(n766), .A2(n764), .ZN(n765) );
  MUX2_X1 U661 ( .A(n4414), .B(DATAIN[31]), .S(n122), .Z(n3497) );
  MUX2_X1 U662 ( .A(n4413), .B(DATAIN[30]), .S(n122), .Z(n3496) );
  MUX2_X1 U663 ( .A(n4412), .B(DATAIN[29]), .S(n122), .Z(n3495) );
  MUX2_X1 U664 ( .A(n4411), .B(DATAIN[28]), .S(n122), .Z(n3494) );
  MUX2_X1 U665 ( .A(n4410), .B(DATAIN[27]), .S(n122), .Z(n3493) );
  MUX2_X1 U666 ( .A(n4409), .B(DATAIN[26]), .S(n122), .Z(n3492) );
  MUX2_X1 U667 ( .A(n4408), .B(DATAIN[25]), .S(n122), .Z(n3491) );
  MUX2_X1 U668 ( .A(n4407), .B(DATAIN[24]), .S(n122), .Z(n3490) );
  MUX2_X1 U669 ( .A(n4406), .B(DATAIN[23]), .S(n121), .Z(n3489) );
  MUX2_X1 U670 ( .A(n4405), .B(DATAIN[22]), .S(n121), .Z(n3488) );
  MUX2_X1 U671 ( .A(n4404), .B(DATAIN[21]), .S(n121), .Z(n3487) );
  MUX2_X1 U672 ( .A(n4403), .B(DATAIN[20]), .S(n121), .Z(n3486) );
  MUX2_X1 U673 ( .A(n4402), .B(DATAIN[19]), .S(n121), .Z(n3485) );
  MUX2_X1 U674 ( .A(n4401), .B(DATAIN[18]), .S(n121), .Z(n3484) );
  MUX2_X1 U675 ( .A(n4400), .B(DATAIN[17]), .S(n121), .Z(n3483) );
  MUX2_X1 U676 ( .A(n4399), .B(DATAIN[16]), .S(n121), .Z(n3482) );
  MUX2_X1 U677 ( .A(n4398), .B(DATAIN[15]), .S(n121), .Z(n3481) );
  MUX2_X1 U678 ( .A(n4397), .B(DATAIN[14]), .S(n121), .Z(n3480) );
  MUX2_X1 U679 ( .A(n4396), .B(DATAIN[13]), .S(n121), .Z(n3479) );
  MUX2_X1 U680 ( .A(n4395), .B(DATAIN[12]), .S(n121), .Z(n3478) );
  MUX2_X1 U681 ( .A(n4394), .B(DATAIN[11]), .S(n120), .Z(n3477) );
  MUX2_X1 U682 ( .A(n4393), .B(DATAIN[10]), .S(n120), .Z(n3476) );
  MUX2_X1 U683 ( .A(n4392), .B(DATAIN[9]), .S(n120), .Z(n3475) );
  MUX2_X1 U684 ( .A(n4391), .B(DATAIN[8]), .S(n120), .Z(n3474) );
  MUX2_X1 U685 ( .A(n4390), .B(DATAIN[7]), .S(n120), .Z(n3473) );
  MUX2_X1 U686 ( .A(n4389), .B(DATAIN[6]), .S(n120), .Z(n3472) );
  MUX2_X1 U687 ( .A(n4388), .B(DATAIN[5]), .S(n120), .Z(n3471) );
  MUX2_X1 U688 ( .A(n4387), .B(DATAIN[4]), .S(n120), .Z(n3470) );
  MUX2_X1 U689 ( .A(n4386), .B(DATAIN[3]), .S(n120), .Z(n3469) );
  MUX2_X1 U690 ( .A(n4385), .B(DATAIN[2]), .S(n120), .Z(n3468) );
  MUX2_X1 U691 ( .A(n4384), .B(DATAIN[1]), .S(n120), .Z(n3467) );
  MUX2_X1 U692 ( .A(n4383), .B(DATAIN[0]), .S(n120), .Z(n3466) );
  AND2_X1 U693 ( .A1(n768), .A2(n764), .ZN(n767) );
  MUX2_X1 U694 ( .A(n769), .B(DATAIN[31]), .S(n125), .Z(n3465) );
  MUX2_X1 U695 ( .A(n771), .B(DATAIN[30]), .S(n125), .Z(n3464) );
  MUX2_X1 U696 ( .A(n772), .B(DATAIN[29]), .S(n125), .Z(n3463) );
  MUX2_X1 U697 ( .A(n773), .B(DATAIN[28]), .S(n125), .Z(n3462) );
  MUX2_X1 U698 ( .A(n774), .B(DATAIN[27]), .S(n125), .Z(n3461) );
  MUX2_X1 U699 ( .A(n775), .B(DATAIN[26]), .S(n125), .Z(n3460) );
  MUX2_X1 U700 ( .A(n776), .B(DATAIN[25]), .S(n125), .Z(n3459) );
  MUX2_X1 U701 ( .A(n777), .B(DATAIN[24]), .S(n125), .Z(n3458) );
  MUX2_X1 U702 ( .A(n778), .B(DATAIN[23]), .S(n124), .Z(n3457) );
  MUX2_X1 U703 ( .A(n779), .B(DATAIN[22]), .S(n124), .Z(n3456) );
  MUX2_X1 U704 ( .A(n780), .B(DATAIN[21]), .S(n124), .Z(n3455) );
  MUX2_X1 U705 ( .A(n781), .B(DATAIN[20]), .S(n124), .Z(n3454) );
  MUX2_X1 U706 ( .A(n782), .B(DATAIN[19]), .S(n124), .Z(n3453) );
  MUX2_X1 U707 ( .A(n783), .B(DATAIN[18]), .S(n124), .Z(n3452) );
  MUX2_X1 U708 ( .A(n784), .B(DATAIN[17]), .S(n124), .Z(n3451) );
  MUX2_X1 U709 ( .A(n785), .B(DATAIN[16]), .S(n124), .Z(n3450) );
  MUX2_X1 U710 ( .A(n786), .B(DATAIN[15]), .S(n124), .Z(n3449) );
  MUX2_X1 U711 ( .A(n787), .B(DATAIN[14]), .S(n124), .Z(n3448) );
  MUX2_X1 U712 ( .A(n788), .B(DATAIN[13]), .S(n124), .Z(n3447) );
  MUX2_X1 U713 ( .A(n789), .B(DATAIN[12]), .S(n124), .Z(n3446) );
  MUX2_X1 U714 ( .A(n790), .B(DATAIN[11]), .S(n123), .Z(n3445) );
  MUX2_X1 U715 ( .A(n791), .B(DATAIN[10]), .S(n123), .Z(n3444) );
  MUX2_X1 U716 ( .A(n792), .B(DATAIN[9]), .S(n123), .Z(n3443) );
  MUX2_X1 U717 ( .A(n793), .B(DATAIN[8]), .S(n123), .Z(n3442) );
  MUX2_X1 U718 ( .A(n794), .B(DATAIN[7]), .S(n123), .Z(n3441) );
  MUX2_X1 U719 ( .A(n795), .B(DATAIN[6]), .S(n123), .Z(n3440) );
  MUX2_X1 U720 ( .A(n796), .B(DATAIN[5]), .S(n123), .Z(n3439) );
  MUX2_X1 U721 ( .A(n797), .B(DATAIN[4]), .S(n123), .Z(n3438) );
  MUX2_X1 U722 ( .A(n798), .B(DATAIN[3]), .S(n123), .Z(n3437) );
  MUX2_X1 U723 ( .A(n799), .B(DATAIN[2]), .S(n123), .Z(n3436) );
  MUX2_X1 U724 ( .A(n800), .B(DATAIN[1]), .S(n123), .Z(n3435) );
  MUX2_X1 U725 ( .A(n801), .B(DATAIN[0]), .S(n123), .Z(n3434) );
  AND2_X1 U726 ( .A1(n802), .A2(n764), .ZN(n770) );
  MUX2_X1 U727 ( .A(n803), .B(DATAIN[31]), .S(n128), .Z(n3433) );
  MUX2_X1 U728 ( .A(n805), .B(DATAIN[30]), .S(n128), .Z(n3432) );
  MUX2_X1 U729 ( .A(n806), .B(DATAIN[29]), .S(n128), .Z(n3431) );
  MUX2_X1 U730 ( .A(n807), .B(DATAIN[28]), .S(n128), .Z(n3430) );
  MUX2_X1 U731 ( .A(n808), .B(DATAIN[27]), .S(n128), .Z(n3429) );
  MUX2_X1 U732 ( .A(n809), .B(DATAIN[26]), .S(n128), .Z(n3428) );
  MUX2_X1 U733 ( .A(n810), .B(DATAIN[25]), .S(n128), .Z(n3427) );
  MUX2_X1 U734 ( .A(n811), .B(DATAIN[24]), .S(n128), .Z(n3426) );
  MUX2_X1 U735 ( .A(n812), .B(DATAIN[23]), .S(n127), .Z(n3425) );
  MUX2_X1 U736 ( .A(n813), .B(DATAIN[22]), .S(n127), .Z(n3424) );
  MUX2_X1 U737 ( .A(n814), .B(DATAIN[21]), .S(n127), .Z(n3423) );
  MUX2_X1 U738 ( .A(n815), .B(DATAIN[20]), .S(n127), .Z(n3422) );
  MUX2_X1 U739 ( .A(n816), .B(DATAIN[19]), .S(n127), .Z(n3421) );
  MUX2_X1 U740 ( .A(n817), .B(DATAIN[18]), .S(n127), .Z(n3420) );
  MUX2_X1 U741 ( .A(n818), .B(DATAIN[17]), .S(n127), .Z(n3419) );
  MUX2_X1 U742 ( .A(n819), .B(DATAIN[16]), .S(n127), .Z(n3418) );
  MUX2_X1 U743 ( .A(n820), .B(DATAIN[15]), .S(n127), .Z(n3417) );
  MUX2_X1 U744 ( .A(n821), .B(DATAIN[14]), .S(n127), .Z(n3416) );
  MUX2_X1 U745 ( .A(n822), .B(DATAIN[13]), .S(n127), .Z(n3415) );
  MUX2_X1 U746 ( .A(n823), .B(DATAIN[12]), .S(n127), .Z(n3414) );
  MUX2_X1 U747 ( .A(n824), .B(DATAIN[11]), .S(n126), .Z(n3413) );
  MUX2_X1 U748 ( .A(n825), .B(DATAIN[10]), .S(n126), .Z(n3412) );
  MUX2_X1 U749 ( .A(n826), .B(DATAIN[9]), .S(n126), .Z(n3411) );
  MUX2_X1 U750 ( .A(n827), .B(DATAIN[8]), .S(n126), .Z(n3410) );
  MUX2_X1 U751 ( .A(n828), .B(DATAIN[7]), .S(n126), .Z(n3409) );
  MUX2_X1 U752 ( .A(n829), .B(DATAIN[6]), .S(n126), .Z(n3408) );
  MUX2_X1 U753 ( .A(n830), .B(DATAIN[5]), .S(n126), .Z(n3407) );
  MUX2_X1 U754 ( .A(n831), .B(DATAIN[4]), .S(n126), .Z(n3406) );
  MUX2_X1 U755 ( .A(n832), .B(DATAIN[3]), .S(n126), .Z(n3405) );
  MUX2_X1 U756 ( .A(n833), .B(DATAIN[2]), .S(n126), .Z(n3404) );
  MUX2_X1 U757 ( .A(n834), .B(DATAIN[1]), .S(n126), .Z(n3403) );
  MUX2_X1 U758 ( .A(n835), .B(DATAIN[0]), .S(n126), .Z(n3402) );
  AND2_X1 U759 ( .A1(n836), .A2(n764), .ZN(n804) );
  MUX2_X1 U760 ( .A(n4382), .B(DATAIN[31]), .S(n131), .Z(n3401) );
  MUX2_X1 U761 ( .A(n4381), .B(DATAIN[30]), .S(n131), .Z(n3400) );
  MUX2_X1 U762 ( .A(n4380), .B(DATAIN[29]), .S(n131), .Z(n3399) );
  MUX2_X1 U763 ( .A(n4379), .B(DATAIN[28]), .S(n131), .Z(n3398) );
  MUX2_X1 U764 ( .A(n4378), .B(DATAIN[27]), .S(n131), .Z(n3397) );
  MUX2_X1 U765 ( .A(n4377), .B(DATAIN[26]), .S(n131), .Z(n3396) );
  MUX2_X1 U766 ( .A(n4376), .B(DATAIN[25]), .S(n131), .Z(n3395) );
  MUX2_X1 U767 ( .A(n4375), .B(DATAIN[24]), .S(n131), .Z(n3394) );
  MUX2_X1 U768 ( .A(n4374), .B(DATAIN[23]), .S(n130), .Z(n3393) );
  MUX2_X1 U769 ( .A(n4373), .B(DATAIN[22]), .S(n130), .Z(n3392) );
  MUX2_X1 U770 ( .A(n4372), .B(DATAIN[21]), .S(n130), .Z(n3391) );
  MUX2_X1 U771 ( .A(n4371), .B(DATAIN[20]), .S(n130), .Z(n3390) );
  MUX2_X1 U772 ( .A(n4370), .B(DATAIN[19]), .S(n130), .Z(n3389) );
  MUX2_X1 U773 ( .A(n4369), .B(DATAIN[18]), .S(n130), .Z(n3388) );
  MUX2_X1 U774 ( .A(n4368), .B(DATAIN[17]), .S(n130), .Z(n3387) );
  MUX2_X1 U775 ( .A(n4367), .B(DATAIN[16]), .S(n130), .Z(n3386) );
  MUX2_X1 U776 ( .A(n4366), .B(DATAIN[15]), .S(n130), .Z(n3385) );
  MUX2_X1 U777 ( .A(n4365), .B(DATAIN[14]), .S(n130), .Z(n3384) );
  MUX2_X1 U778 ( .A(n4364), .B(DATAIN[13]), .S(n130), .Z(n3383) );
  MUX2_X1 U779 ( .A(n4363), .B(DATAIN[12]), .S(n130), .Z(n3382) );
  MUX2_X1 U780 ( .A(n4362), .B(DATAIN[11]), .S(n129), .Z(n3381) );
  MUX2_X1 U781 ( .A(n4361), .B(DATAIN[10]), .S(n129), .Z(n3380) );
  MUX2_X1 U782 ( .A(n4360), .B(DATAIN[9]), .S(n129), .Z(n3379) );
  MUX2_X1 U783 ( .A(n4359), .B(DATAIN[8]), .S(n129), .Z(n3378) );
  MUX2_X1 U784 ( .A(n4358), .B(DATAIN[7]), .S(n129), .Z(n3377) );
  MUX2_X1 U785 ( .A(n4357), .B(DATAIN[6]), .S(n129), .Z(n3376) );
  MUX2_X1 U786 ( .A(n4356), .B(DATAIN[5]), .S(n129), .Z(n3375) );
  MUX2_X1 U787 ( .A(n4355), .B(DATAIN[4]), .S(n129), .Z(n3374) );
  MUX2_X1 U788 ( .A(n4354), .B(DATAIN[3]), .S(n129), .Z(n3373) );
  MUX2_X1 U789 ( .A(n4353), .B(DATAIN[2]), .S(n129), .Z(n3372) );
  MUX2_X1 U790 ( .A(n4352), .B(DATAIN[1]), .S(n129), .Z(n3371) );
  MUX2_X1 U791 ( .A(n4351), .B(DATAIN[0]), .S(n129), .Z(n3370) );
  AND2_X1 U792 ( .A1(n870), .A2(n764), .ZN(n869) );
  MUX2_X1 U793 ( .A(n4350), .B(DATAIN[31]), .S(n134), .Z(n3369) );
  MUX2_X1 U794 ( .A(n4349), .B(DATAIN[30]), .S(n134), .Z(n3368) );
  MUX2_X1 U795 ( .A(n4348), .B(DATAIN[29]), .S(n134), .Z(n3367) );
  MUX2_X1 U796 ( .A(n4347), .B(DATAIN[28]), .S(n134), .Z(n3366) );
  MUX2_X1 U797 ( .A(n4346), .B(DATAIN[27]), .S(n134), .Z(n3365) );
  MUX2_X1 U798 ( .A(n4345), .B(DATAIN[26]), .S(n134), .Z(n3364) );
  MUX2_X1 U799 ( .A(n4344), .B(DATAIN[25]), .S(n134), .Z(n3363) );
  MUX2_X1 U800 ( .A(n4343), .B(DATAIN[24]), .S(n134), .Z(n3362) );
  MUX2_X1 U801 ( .A(n4342), .B(DATAIN[23]), .S(n133), .Z(n3361) );
  MUX2_X1 U802 ( .A(n4341), .B(DATAIN[22]), .S(n133), .Z(n3360) );
  MUX2_X1 U803 ( .A(n4340), .B(DATAIN[21]), .S(n133), .Z(n3359) );
  MUX2_X1 U804 ( .A(n4339), .B(DATAIN[20]), .S(n133), .Z(n3358) );
  MUX2_X1 U805 ( .A(n4338), .B(DATAIN[19]), .S(n133), .Z(n3357) );
  MUX2_X1 U806 ( .A(n4337), .B(DATAIN[18]), .S(n133), .Z(n3356) );
  MUX2_X1 U807 ( .A(n4336), .B(DATAIN[17]), .S(n133), .Z(n3355) );
  MUX2_X1 U808 ( .A(n4335), .B(DATAIN[16]), .S(n133), .Z(n3354) );
  MUX2_X1 U809 ( .A(n4334), .B(DATAIN[15]), .S(n133), .Z(n3353) );
  MUX2_X1 U810 ( .A(n4333), .B(DATAIN[14]), .S(n133), .Z(n3352) );
  MUX2_X1 U811 ( .A(n4332), .B(DATAIN[13]), .S(n133), .Z(n3351) );
  MUX2_X1 U812 ( .A(n4331), .B(DATAIN[12]), .S(n133), .Z(n3350) );
  MUX2_X1 U813 ( .A(n4330), .B(DATAIN[11]), .S(n132), .Z(n3349) );
  MUX2_X1 U814 ( .A(n4329), .B(DATAIN[10]), .S(n132), .Z(n3348) );
  MUX2_X1 U815 ( .A(n4328), .B(DATAIN[9]), .S(n132), .Z(n3347) );
  MUX2_X1 U816 ( .A(n4327), .B(DATAIN[8]), .S(n132), .Z(n3346) );
  MUX2_X1 U817 ( .A(n4326), .B(DATAIN[7]), .S(n132), .Z(n3345) );
  MUX2_X1 U818 ( .A(n4325), .B(DATAIN[6]), .S(n132), .Z(n3344) );
  MUX2_X1 U819 ( .A(n4324), .B(DATAIN[5]), .S(n132), .Z(n3343) );
  MUX2_X1 U820 ( .A(n4323), .B(DATAIN[4]), .S(n132), .Z(n3342) );
  MUX2_X1 U821 ( .A(n4322), .B(DATAIN[3]), .S(n132), .Z(n3341) );
  MUX2_X1 U822 ( .A(n4321), .B(DATAIN[2]), .S(n132), .Z(n3340) );
  MUX2_X1 U823 ( .A(n4320), .B(DATAIN[1]), .S(n132), .Z(n3339) );
  MUX2_X1 U824 ( .A(n4319), .B(DATAIN[0]), .S(n132), .Z(n3338) );
  AND2_X1 U825 ( .A1(n872), .A2(n764), .ZN(n871) );
  AND3_X1 U826 ( .A1(n873), .A2(n874), .A3(n875), .ZN(n764) );
  INV_X1 U827 ( .A(n876), .ZN(n3337) );
  MUX2_X1 U828 ( .A(n229), .B(n593), .S(n137), .Z(n876) );
  INV_X1 U829 ( .A(n878), .ZN(n3336) );
  MUX2_X1 U830 ( .A(n230), .B(n592), .S(n137), .Z(n878) );
  INV_X1 U831 ( .A(n879), .ZN(n3335) );
  MUX2_X1 U832 ( .A(n231), .B(n591), .S(n137), .Z(n879) );
  INV_X1 U833 ( .A(n880), .ZN(n3334) );
  MUX2_X1 U834 ( .A(n232), .B(n590), .S(n137), .Z(n880) );
  INV_X1 U835 ( .A(n881), .ZN(n3333) );
  MUX2_X1 U836 ( .A(n233), .B(n589), .S(n137), .Z(n881) );
  INV_X1 U837 ( .A(n882), .ZN(n3332) );
  MUX2_X1 U838 ( .A(n234), .B(n588), .S(n137), .Z(n882) );
  INV_X1 U839 ( .A(n883), .ZN(n3331) );
  MUX2_X1 U840 ( .A(n235), .B(n587), .S(n137), .Z(n883) );
  INV_X1 U841 ( .A(n884), .ZN(n3330) );
  MUX2_X1 U842 ( .A(n236), .B(n586), .S(n137), .Z(n884) );
  INV_X1 U843 ( .A(n885), .ZN(n3329) );
  MUX2_X1 U844 ( .A(n237), .B(n585), .S(n136), .Z(n885) );
  INV_X1 U845 ( .A(n886), .ZN(n3328) );
  MUX2_X1 U846 ( .A(n238), .B(n584), .S(n136), .Z(n886) );
  INV_X1 U847 ( .A(n887), .ZN(n3327) );
  MUX2_X1 U848 ( .A(n239), .B(n583), .S(n136), .Z(n887) );
  INV_X1 U849 ( .A(n888), .ZN(n3326) );
  MUX2_X1 U850 ( .A(n240), .B(n582), .S(n136), .Z(n888) );
  INV_X1 U851 ( .A(n889), .ZN(n3325) );
  MUX2_X1 U852 ( .A(n241), .B(n581), .S(n136), .Z(n889) );
  INV_X1 U853 ( .A(n890), .ZN(n3324) );
  MUX2_X1 U854 ( .A(n242), .B(n580), .S(n136), .Z(n890) );
  INV_X1 U855 ( .A(n891), .ZN(n3323) );
  MUX2_X1 U856 ( .A(n243), .B(n579), .S(n136), .Z(n891) );
  INV_X1 U857 ( .A(n892), .ZN(n3322) );
  MUX2_X1 U858 ( .A(n244), .B(n578), .S(n136), .Z(n892) );
  INV_X1 U859 ( .A(n893), .ZN(n3321) );
  MUX2_X1 U860 ( .A(n245), .B(n577), .S(n136), .Z(n893) );
  INV_X1 U861 ( .A(n894), .ZN(n3320) );
  MUX2_X1 U862 ( .A(n246), .B(n576), .S(n136), .Z(n894) );
  INV_X1 U863 ( .A(n895), .ZN(n3319) );
  MUX2_X1 U864 ( .A(n247), .B(n575), .S(n136), .Z(n895) );
  INV_X1 U865 ( .A(n896), .ZN(n3318) );
  MUX2_X1 U866 ( .A(n248), .B(n574), .S(n136), .Z(n896) );
  INV_X1 U867 ( .A(n897), .ZN(n3317) );
  MUX2_X1 U868 ( .A(n249), .B(n573), .S(n135), .Z(n897) );
  INV_X1 U869 ( .A(n898), .ZN(n3316) );
  MUX2_X1 U870 ( .A(n250), .B(n572), .S(n135), .Z(n898) );
  INV_X1 U871 ( .A(n899), .ZN(n3315) );
  MUX2_X1 U872 ( .A(n251), .B(n571), .S(n135), .Z(n899) );
  INV_X1 U873 ( .A(n900), .ZN(n3314) );
  MUX2_X1 U874 ( .A(n252), .B(n570), .S(n135), .Z(n900) );
  INV_X1 U875 ( .A(n901), .ZN(n3313) );
  MUX2_X1 U876 ( .A(n253), .B(n569), .S(n135), .Z(n901) );
  INV_X1 U877 ( .A(n902), .ZN(n3312) );
  MUX2_X1 U878 ( .A(n254), .B(n568), .S(n135), .Z(n902) );
  INV_X1 U879 ( .A(n903), .ZN(n3311) );
  MUX2_X1 U880 ( .A(n255), .B(n567), .S(n135), .Z(n903) );
  INV_X1 U881 ( .A(n904), .ZN(n3310) );
  MUX2_X1 U882 ( .A(n256), .B(n566), .S(n135), .Z(n904) );
  INV_X1 U883 ( .A(n905), .ZN(n3309) );
  MUX2_X1 U884 ( .A(n257), .B(n565), .S(n135), .Z(n905) );
  INV_X1 U885 ( .A(n906), .ZN(n3308) );
  MUX2_X1 U886 ( .A(n258), .B(n564), .S(n135), .Z(n906) );
  INV_X1 U887 ( .A(n907), .ZN(n3307) );
  MUX2_X1 U888 ( .A(n259), .B(n563), .S(n135), .Z(n907) );
  INV_X1 U889 ( .A(n908), .ZN(n3306) );
  MUX2_X1 U890 ( .A(n260), .B(n562), .S(n135), .Z(n908) );
  AND2_X1 U891 ( .A1(n909), .A2(n910), .ZN(n877) );
  INV_X1 U892 ( .A(n911), .ZN(n3305) );
  MUX2_X1 U893 ( .A(n261), .B(n593), .S(n140), .Z(n911) );
  INV_X1 U894 ( .A(n913), .ZN(n3304) );
  MUX2_X1 U895 ( .A(n262), .B(n592), .S(n140), .Z(n913) );
  INV_X1 U896 ( .A(n914), .ZN(n3303) );
  MUX2_X1 U897 ( .A(n263), .B(n591), .S(n140), .Z(n914) );
  INV_X1 U898 ( .A(n915), .ZN(n3302) );
  MUX2_X1 U899 ( .A(n264), .B(n590), .S(n140), .Z(n915) );
  INV_X1 U900 ( .A(n916), .ZN(n3301) );
  MUX2_X1 U901 ( .A(n265), .B(n589), .S(n140), .Z(n916) );
  INV_X1 U902 ( .A(n917), .ZN(n3300) );
  MUX2_X1 U903 ( .A(n266), .B(n588), .S(n140), .Z(n917) );
  INV_X1 U904 ( .A(n918), .ZN(n3299) );
  MUX2_X1 U905 ( .A(n267), .B(n587), .S(n140), .Z(n918) );
  INV_X1 U906 ( .A(n919), .ZN(n3298) );
  MUX2_X1 U907 ( .A(n268), .B(n586), .S(n140), .Z(n919) );
  INV_X1 U908 ( .A(n920), .ZN(n3297) );
  MUX2_X1 U909 ( .A(n269), .B(n585), .S(n139), .Z(n920) );
  INV_X1 U910 ( .A(n921), .ZN(n3296) );
  MUX2_X1 U911 ( .A(n270), .B(n584), .S(n139), .Z(n921) );
  INV_X1 U912 ( .A(n922), .ZN(n3295) );
  MUX2_X1 U913 ( .A(n271), .B(n583), .S(n139), .Z(n922) );
  INV_X1 U914 ( .A(n923), .ZN(n3294) );
  MUX2_X1 U915 ( .A(n272), .B(n582), .S(n139), .Z(n923) );
  INV_X1 U916 ( .A(n924), .ZN(n3293) );
  MUX2_X1 U917 ( .A(n273), .B(n581), .S(n139), .Z(n924) );
  INV_X1 U918 ( .A(n925), .ZN(n3292) );
  MUX2_X1 U919 ( .A(n274), .B(n580), .S(n139), .Z(n925) );
  INV_X1 U920 ( .A(n926), .ZN(n3291) );
  MUX2_X1 U921 ( .A(n275), .B(n579), .S(n139), .Z(n926) );
  INV_X1 U922 ( .A(n927), .ZN(n3290) );
  MUX2_X1 U923 ( .A(n276), .B(n578), .S(n139), .Z(n927) );
  INV_X1 U924 ( .A(n928), .ZN(n3289) );
  MUX2_X1 U925 ( .A(n277), .B(n577), .S(n139), .Z(n928) );
  INV_X1 U926 ( .A(n929), .ZN(n3288) );
  MUX2_X1 U927 ( .A(n278), .B(n576), .S(n139), .Z(n929) );
  INV_X1 U928 ( .A(n930), .ZN(n3287) );
  MUX2_X1 U929 ( .A(n279), .B(n575), .S(n139), .Z(n930) );
  INV_X1 U930 ( .A(n931), .ZN(n3286) );
  MUX2_X1 U931 ( .A(n280), .B(n574), .S(n139), .Z(n931) );
  INV_X1 U932 ( .A(n932), .ZN(n3285) );
  MUX2_X1 U933 ( .A(n281), .B(n573), .S(n138), .Z(n932) );
  INV_X1 U934 ( .A(n965), .ZN(n3284) );
  MUX2_X1 U935 ( .A(n282), .B(n572), .S(n138), .Z(n965) );
  INV_X1 U936 ( .A(n966), .ZN(n3283) );
  MUX2_X1 U937 ( .A(n283), .B(n571), .S(n138), .Z(n966) );
  INV_X1 U938 ( .A(n967), .ZN(n3282) );
  MUX2_X1 U939 ( .A(n284), .B(n570), .S(n138), .Z(n967) );
  INV_X1 U940 ( .A(n968), .ZN(n3281) );
  MUX2_X1 U941 ( .A(n285), .B(n569), .S(n138), .Z(n968) );
  INV_X1 U942 ( .A(n969), .ZN(n3280) );
  MUX2_X1 U943 ( .A(n286), .B(n568), .S(n138), .Z(n969) );
  INV_X1 U944 ( .A(n970), .ZN(n3279) );
  MUX2_X1 U945 ( .A(n287), .B(n567), .S(n138), .Z(n970) );
  INV_X1 U946 ( .A(n971), .ZN(n3278) );
  MUX2_X1 U947 ( .A(n288), .B(n566), .S(n138), .Z(n971) );
  INV_X1 U948 ( .A(n972), .ZN(n3277) );
  MUX2_X1 U949 ( .A(n289), .B(n565), .S(n138), .Z(n972) );
  INV_X1 U950 ( .A(n973), .ZN(n3276) );
  MUX2_X1 U951 ( .A(n290), .B(n564), .S(n138), .Z(n973) );
  INV_X1 U952 ( .A(n974), .ZN(n3275) );
  MUX2_X1 U953 ( .A(n291), .B(n563), .S(n138), .Z(n974) );
  INV_X1 U954 ( .A(n975), .ZN(n3274) );
  MUX2_X1 U955 ( .A(n292), .B(n562), .S(n138), .Z(n975) );
  AND2_X1 U956 ( .A1(n909), .A2(n763), .ZN(n912) );
  MUX2_X1 U957 ( .A(n4318), .B(DATAIN[31]), .S(n143), .Z(n3273) );
  MUX2_X1 U958 ( .A(n4317), .B(DATAIN[30]), .S(n143), .Z(n3272) );
  MUX2_X1 U959 ( .A(n4316), .B(DATAIN[29]), .S(n143), .Z(n3271) );
  MUX2_X1 U960 ( .A(n4315), .B(DATAIN[28]), .S(n143), .Z(n3270) );
  MUX2_X1 U961 ( .A(n4314), .B(DATAIN[27]), .S(n143), .Z(n3269) );
  MUX2_X1 U962 ( .A(n4313), .B(DATAIN[26]), .S(n143), .Z(n3268) );
  MUX2_X1 U963 ( .A(n4312), .B(DATAIN[25]), .S(n143), .Z(n3267) );
  MUX2_X1 U964 ( .A(n4311), .B(DATAIN[24]), .S(n143), .Z(n3266) );
  MUX2_X1 U965 ( .A(n4310), .B(DATAIN[23]), .S(n142), .Z(n3265) );
  MUX2_X1 U966 ( .A(n4309), .B(DATAIN[22]), .S(n142), .Z(n3264) );
  MUX2_X1 U967 ( .A(n4308), .B(DATAIN[21]), .S(n142), .Z(n3263) );
  MUX2_X1 U968 ( .A(n4307), .B(DATAIN[20]), .S(n142), .Z(n3262) );
  MUX2_X1 U969 ( .A(n4306), .B(DATAIN[19]), .S(n142), .Z(n3261) );
  MUX2_X1 U970 ( .A(n4305), .B(DATAIN[18]), .S(n142), .Z(n3260) );
  MUX2_X1 U971 ( .A(n4304), .B(DATAIN[17]), .S(n142), .Z(n3259) );
  MUX2_X1 U972 ( .A(n4303), .B(DATAIN[16]), .S(n142), .Z(n3258) );
  MUX2_X1 U973 ( .A(n4302), .B(DATAIN[15]), .S(n142), .Z(n3257) );
  MUX2_X1 U974 ( .A(n4301), .B(DATAIN[14]), .S(n142), .Z(n3256) );
  MUX2_X1 U975 ( .A(n4300), .B(DATAIN[13]), .S(n142), .Z(n3255) );
  MUX2_X1 U976 ( .A(n4299), .B(DATAIN[12]), .S(n142), .Z(n3254) );
  MUX2_X1 U977 ( .A(n4298), .B(DATAIN[11]), .S(n141), .Z(n3253) );
  MUX2_X1 U978 ( .A(n4297), .B(DATAIN[10]), .S(n141), .Z(n3252) );
  MUX2_X1 U979 ( .A(n4296), .B(DATAIN[9]), .S(n141), .Z(n3251) );
  MUX2_X1 U980 ( .A(n4295), .B(DATAIN[8]), .S(n141), .Z(n3250) );
  MUX2_X1 U981 ( .A(n4294), .B(DATAIN[7]), .S(n141), .Z(n3249) );
  MUX2_X1 U982 ( .A(n4293), .B(DATAIN[6]), .S(n141), .Z(n3248) );
  MUX2_X1 U983 ( .A(n4292), .B(DATAIN[5]), .S(n141), .Z(n3247) );
  MUX2_X1 U984 ( .A(n4291), .B(DATAIN[4]), .S(n141), .Z(n3246) );
  MUX2_X1 U985 ( .A(n4290), .B(DATAIN[3]), .S(n141), .Z(n3245) );
  MUX2_X1 U986 ( .A(n4289), .B(DATAIN[2]), .S(n141), .Z(n3244) );
  MUX2_X1 U987 ( .A(n4288), .B(DATAIN[1]), .S(n141), .Z(n3243) );
  MUX2_X1 U988 ( .A(n4287), .B(DATAIN[0]), .S(n141), .Z(n3242) );
  AND2_X1 U989 ( .A1(n909), .A2(n766), .ZN(n976) );
  MUX2_X1 U990 ( .A(n4286), .B(DATAIN[31]), .S(n146), .Z(n3241) );
  MUX2_X1 U991 ( .A(n4285), .B(DATAIN[30]), .S(n146), .Z(n3240) );
  MUX2_X1 U992 ( .A(n4284), .B(DATAIN[29]), .S(n146), .Z(n3239) );
  MUX2_X1 U993 ( .A(n4283), .B(DATAIN[28]), .S(n146), .Z(n3238) );
  MUX2_X1 U994 ( .A(n4282), .B(DATAIN[27]), .S(n146), .Z(n3237) );
  MUX2_X1 U995 ( .A(n4281), .B(DATAIN[26]), .S(n146), .Z(n3236) );
  MUX2_X1 U996 ( .A(n4280), .B(DATAIN[25]), .S(n146), .Z(n3235) );
  MUX2_X1 U997 ( .A(n4279), .B(DATAIN[24]), .S(n146), .Z(n3234) );
  MUX2_X1 U998 ( .A(n4278), .B(DATAIN[23]), .S(n145), .Z(n3233) );
  MUX2_X1 U999 ( .A(n4277), .B(DATAIN[22]), .S(n145), .Z(n3232) );
  MUX2_X1 U1000 ( .A(n4276), .B(DATAIN[21]), .S(n145), .Z(n3231) );
  MUX2_X1 U1001 ( .A(n4275), .B(DATAIN[20]), .S(n145), .Z(n3230) );
  MUX2_X1 U1002 ( .A(n4274), .B(DATAIN[19]), .S(n145), .Z(n3229) );
  MUX2_X1 U1003 ( .A(n4273), .B(DATAIN[18]), .S(n145), .Z(n3228) );
  MUX2_X1 U1004 ( .A(n4272), .B(DATAIN[17]), .S(n145), .Z(n3227) );
  MUX2_X1 U1005 ( .A(n4271), .B(DATAIN[16]), .S(n145), .Z(n3226) );
  MUX2_X1 U1006 ( .A(n4270), .B(DATAIN[15]), .S(n145), .Z(n3225) );
  MUX2_X1 U1007 ( .A(n4269), .B(DATAIN[14]), .S(n145), .Z(n3224) );
  MUX2_X1 U1008 ( .A(n4268), .B(DATAIN[13]), .S(n145), .Z(n3223) );
  MUX2_X1 U1009 ( .A(n4267), .B(DATAIN[12]), .S(n145), .Z(n3222) );
  MUX2_X1 U1010 ( .A(n4266), .B(DATAIN[11]), .S(n144), .Z(n3221) );
  MUX2_X1 U1011 ( .A(n4265), .B(DATAIN[10]), .S(n144), .Z(n3220) );
  MUX2_X1 U1012 ( .A(n4264), .B(DATAIN[9]), .S(n144), .Z(n3219) );
  MUX2_X1 U1013 ( .A(n4263), .B(DATAIN[8]), .S(n144), .Z(n3218) );
  MUX2_X1 U1014 ( .A(n4262), .B(DATAIN[7]), .S(n144), .Z(n3217) );
  MUX2_X1 U1015 ( .A(n4261), .B(DATAIN[6]), .S(n144), .Z(n3216) );
  MUX2_X1 U1016 ( .A(n4260), .B(DATAIN[5]), .S(n144), .Z(n3215) );
  MUX2_X1 U1017 ( .A(n4259), .B(DATAIN[4]), .S(n144), .Z(n3214) );
  MUX2_X1 U1018 ( .A(n4258), .B(DATAIN[3]), .S(n144), .Z(n3213) );
  MUX2_X1 U1019 ( .A(n4257), .B(DATAIN[2]), .S(n144), .Z(n3212) );
  MUX2_X1 U1020 ( .A(n4256), .B(DATAIN[1]), .S(n144), .Z(n3211) );
  MUX2_X1 U1021 ( .A(n4255), .B(DATAIN[0]), .S(n144), .Z(n3210) );
  AND2_X1 U1022 ( .A1(n909), .A2(n768), .ZN(n977) );
  INV_X1 U1023 ( .A(n978), .ZN(n3209) );
  MUX2_X1 U1024 ( .A(n357), .B(n593), .S(n149), .Z(n978) );
  INV_X1 U1025 ( .A(n980), .ZN(n3208) );
  MUX2_X1 U1026 ( .A(n358), .B(n592), .S(n149), .Z(n980) );
  INV_X1 U1027 ( .A(n981), .ZN(n3207) );
  MUX2_X1 U1028 ( .A(n359), .B(n591), .S(n149), .Z(n981) );
  INV_X1 U1029 ( .A(n982), .ZN(n3206) );
  MUX2_X1 U1030 ( .A(n360), .B(n590), .S(n149), .Z(n982) );
  INV_X1 U1031 ( .A(n983), .ZN(n3205) );
  MUX2_X1 U1032 ( .A(n361), .B(n589), .S(n149), .Z(n983) );
  INV_X1 U1033 ( .A(n984), .ZN(n3204) );
  MUX2_X1 U1034 ( .A(n362), .B(n588), .S(n149), .Z(n984) );
  INV_X1 U1035 ( .A(n985), .ZN(n3203) );
  MUX2_X1 U1036 ( .A(n363), .B(n587), .S(n149), .Z(n985) );
  INV_X1 U1037 ( .A(n986), .ZN(n3202) );
  MUX2_X1 U1038 ( .A(n364), .B(n586), .S(n149), .Z(n986) );
  INV_X1 U1039 ( .A(n987), .ZN(n3201) );
  MUX2_X1 U1040 ( .A(n365), .B(n585), .S(n148), .Z(n987) );
  INV_X1 U1041 ( .A(n988), .ZN(n3200) );
  MUX2_X1 U1042 ( .A(n366), .B(n584), .S(n148), .Z(n988) );
  INV_X1 U1043 ( .A(n989), .ZN(n3199) );
  MUX2_X1 U1044 ( .A(n367), .B(n583), .S(n148), .Z(n989) );
  INV_X1 U1045 ( .A(n990), .ZN(n3198) );
  MUX2_X1 U1046 ( .A(n368), .B(n582), .S(n148), .Z(n990) );
  INV_X1 U1047 ( .A(n991), .ZN(n3197) );
  MUX2_X1 U1048 ( .A(n369), .B(n581), .S(n148), .Z(n991) );
  INV_X1 U1049 ( .A(n992), .ZN(n3196) );
  MUX2_X1 U1050 ( .A(n370), .B(n580), .S(n148), .Z(n992) );
  INV_X1 U1051 ( .A(n993), .ZN(n3195) );
  MUX2_X1 U1052 ( .A(n371), .B(n579), .S(n148), .Z(n993) );
  INV_X1 U1053 ( .A(n994), .ZN(n3194) );
  MUX2_X1 U1054 ( .A(n372), .B(n578), .S(n148), .Z(n994) );
  INV_X1 U1055 ( .A(n995), .ZN(n3193) );
  MUX2_X1 U1056 ( .A(n373), .B(n577), .S(n148), .Z(n995) );
  INV_X1 U1057 ( .A(n996), .ZN(n3192) );
  MUX2_X1 U1058 ( .A(n374), .B(n576), .S(n148), .Z(n996) );
  INV_X1 U1059 ( .A(n997), .ZN(n3191) );
  MUX2_X1 U1060 ( .A(n375), .B(n575), .S(n148), .Z(n997) );
  INV_X1 U1061 ( .A(n998), .ZN(n3190) );
  MUX2_X1 U1062 ( .A(n376), .B(n574), .S(n148), .Z(n998) );
  INV_X1 U1063 ( .A(n999), .ZN(n3189) );
  MUX2_X1 U1064 ( .A(n377), .B(n573), .S(n147), .Z(n999) );
  INV_X1 U1065 ( .A(n1000), .ZN(n3188) );
  MUX2_X1 U1066 ( .A(n378), .B(n572), .S(n147), .Z(n1000) );
  INV_X1 U1067 ( .A(n1001), .ZN(n3187) );
  MUX2_X1 U1068 ( .A(n379), .B(n571), .S(n147), .Z(n1001) );
  INV_X1 U1069 ( .A(n1002), .ZN(n3186) );
  MUX2_X1 U1070 ( .A(n380), .B(n570), .S(n147), .Z(n1002) );
  INV_X1 U1071 ( .A(n1003), .ZN(n3185) );
  MUX2_X1 U1072 ( .A(n381), .B(n569), .S(n147), .Z(n1003) );
  INV_X1 U1073 ( .A(n1004), .ZN(n3184) );
  MUX2_X1 U1074 ( .A(n382), .B(n568), .S(n147), .Z(n1004) );
  INV_X1 U1075 ( .A(n1005), .ZN(n3183) );
  MUX2_X1 U1076 ( .A(n383), .B(n567), .S(n147), .Z(n1005) );
  INV_X1 U1077 ( .A(n1006), .ZN(n3182) );
  MUX2_X1 U1078 ( .A(n384), .B(n566), .S(n147), .Z(n1006) );
  INV_X1 U1079 ( .A(n1007), .ZN(n3181) );
  MUX2_X1 U1080 ( .A(n385), .B(n565), .S(n147), .Z(n1007) );
  INV_X1 U1081 ( .A(n1008), .ZN(n3180) );
  MUX2_X1 U1082 ( .A(n386), .B(n564), .S(n147), .Z(n1008) );
  INV_X1 U1083 ( .A(n1009), .ZN(n3179) );
  MUX2_X1 U1084 ( .A(n387), .B(n563), .S(n147), .Z(n1009) );
  INV_X1 U1085 ( .A(n1010), .ZN(n3178) );
  MUX2_X1 U1086 ( .A(n388), .B(n562), .S(n147), .Z(n1010) );
  AND2_X1 U1087 ( .A1(n909), .A2(n802), .ZN(n979) );
  INV_X1 U1088 ( .A(n1011), .ZN(n3177) );
  MUX2_X1 U1089 ( .A(n389), .B(n593), .S(n152), .Z(n1011) );
  INV_X1 U1090 ( .A(n1013), .ZN(n3176) );
  MUX2_X1 U1091 ( .A(n390), .B(n592), .S(n152), .Z(n1013) );
  INV_X1 U1092 ( .A(n1014), .ZN(n3175) );
  MUX2_X1 U1093 ( .A(n391), .B(n591), .S(n152), .Z(n1014) );
  INV_X1 U1094 ( .A(n1015), .ZN(n3174) );
  MUX2_X1 U1095 ( .A(n392), .B(n590), .S(n152), .Z(n1015) );
  INV_X1 U1096 ( .A(n1016), .ZN(n3173) );
  MUX2_X1 U1097 ( .A(n393), .B(n589), .S(n152), .Z(n1016) );
  INV_X1 U1098 ( .A(n1017), .ZN(n3172) );
  MUX2_X1 U1099 ( .A(n394), .B(n588), .S(n152), .Z(n1017) );
  INV_X1 U1100 ( .A(n1018), .ZN(n3171) );
  MUX2_X1 U1101 ( .A(n395), .B(n587), .S(n152), .Z(n1018) );
  INV_X1 U1102 ( .A(n1019), .ZN(n3170) );
  MUX2_X1 U1103 ( .A(n396), .B(n586), .S(n152), .Z(n1019) );
  INV_X1 U1104 ( .A(n1020), .ZN(n3169) );
  MUX2_X1 U1105 ( .A(n397), .B(n585), .S(n151), .Z(n1020) );
  INV_X1 U1106 ( .A(n1021), .ZN(n3168) );
  MUX2_X1 U1107 ( .A(n398), .B(n584), .S(n151), .Z(n1021) );
  INV_X1 U1108 ( .A(n1022), .ZN(n3167) );
  MUX2_X1 U1109 ( .A(n399), .B(n583), .S(n151), .Z(n1022) );
  INV_X1 U1110 ( .A(n1023), .ZN(n3166) );
  MUX2_X1 U1111 ( .A(n400), .B(n582), .S(n151), .Z(n1023) );
  INV_X1 U1112 ( .A(n1024), .ZN(n3165) );
  MUX2_X1 U1113 ( .A(n401), .B(n581), .S(n151), .Z(n1024) );
  INV_X1 U1114 ( .A(n1025), .ZN(n3164) );
  MUX2_X1 U1115 ( .A(n402), .B(n580), .S(n151), .Z(n1025) );
  INV_X1 U1116 ( .A(n1026), .ZN(n3163) );
  MUX2_X1 U1117 ( .A(n403), .B(n579), .S(n151), .Z(n1026) );
  INV_X1 U1118 ( .A(n1027), .ZN(n3162) );
  MUX2_X1 U1119 ( .A(n404), .B(n578), .S(n151), .Z(n1027) );
  INV_X1 U1120 ( .A(n1028), .ZN(n3161) );
  MUX2_X1 U1121 ( .A(n405), .B(n577), .S(n151), .Z(n1028) );
  INV_X1 U1122 ( .A(n1029), .ZN(n3160) );
  MUX2_X1 U1123 ( .A(n406), .B(n576), .S(n151), .Z(n1029) );
  INV_X1 U1124 ( .A(n1030), .ZN(n3159) );
  MUX2_X1 U1125 ( .A(n407), .B(n575), .S(n151), .Z(n1030) );
  INV_X1 U1126 ( .A(n1031), .ZN(n3158) );
  MUX2_X1 U1127 ( .A(n408), .B(n574), .S(n151), .Z(n1031) );
  INV_X1 U1128 ( .A(n1032), .ZN(n3157) );
  MUX2_X1 U1129 ( .A(n409), .B(n573), .S(n150), .Z(n1032) );
  INV_X1 U1130 ( .A(n1033), .ZN(n3156) );
  MUX2_X1 U1131 ( .A(n410), .B(n572), .S(n150), .Z(n1033) );
  INV_X1 U1132 ( .A(n1034), .ZN(n3155) );
  MUX2_X1 U1133 ( .A(n411), .B(n571), .S(n150), .Z(n1034) );
  INV_X1 U1134 ( .A(n1035), .ZN(n3154) );
  MUX2_X1 U1135 ( .A(n412), .B(n570), .S(n150), .Z(n1035) );
  INV_X1 U1136 ( .A(n1036), .ZN(n3153) );
  MUX2_X1 U1137 ( .A(n413), .B(n569), .S(n150), .Z(n1036) );
  INV_X1 U1138 ( .A(n1037), .ZN(n3152) );
  MUX2_X1 U1139 ( .A(n414), .B(n568), .S(n150), .Z(n1037) );
  INV_X1 U1140 ( .A(n1038), .ZN(n3151) );
  MUX2_X1 U1141 ( .A(n415), .B(n567), .S(n150), .Z(n1038) );
  INV_X1 U1142 ( .A(n1039), .ZN(n3150) );
  MUX2_X1 U1143 ( .A(n416), .B(n566), .S(n150), .Z(n1039) );
  INV_X1 U1144 ( .A(n1040), .ZN(n3149) );
  MUX2_X1 U1145 ( .A(n417), .B(n565), .S(n150), .Z(n1040) );
  INV_X1 U1146 ( .A(n1041), .ZN(n3148) );
  MUX2_X1 U1147 ( .A(n418), .B(n564), .S(n150), .Z(n1041) );
  INV_X1 U1148 ( .A(n1042), .ZN(n3147) );
  MUX2_X1 U1149 ( .A(n419), .B(n563), .S(n150), .Z(n1042) );
  INV_X1 U1150 ( .A(n1043), .ZN(n3146) );
  MUX2_X1 U1151 ( .A(n420), .B(n562), .S(n150), .Z(n1043) );
  AND2_X1 U1152 ( .A1(n909), .A2(n836), .ZN(n1012) );
  MUX2_X1 U1153 ( .A(n4254), .B(DATAIN[31]), .S(n155), .Z(n3145) );
  MUX2_X1 U1154 ( .A(n4253), .B(DATAIN[30]), .S(n155), .Z(n3144) );
  MUX2_X1 U1155 ( .A(n4252), .B(DATAIN[29]), .S(n155), .Z(n3143) );
  MUX2_X1 U1156 ( .A(n4251), .B(DATAIN[28]), .S(n155), .Z(n3142) );
  MUX2_X1 U1157 ( .A(n4250), .B(DATAIN[27]), .S(n155), .Z(n3141) );
  MUX2_X1 U1158 ( .A(n4249), .B(DATAIN[26]), .S(n155), .Z(n3140) );
  MUX2_X1 U1159 ( .A(n4248), .B(DATAIN[25]), .S(n155), .Z(n3139) );
  MUX2_X1 U1160 ( .A(n4247), .B(DATAIN[24]), .S(n155), .Z(n3138) );
  MUX2_X1 U1161 ( .A(n4246), .B(DATAIN[23]), .S(n154), .Z(n3137) );
  MUX2_X1 U1162 ( .A(n4245), .B(DATAIN[22]), .S(n154), .Z(n3136) );
  MUX2_X1 U1163 ( .A(n4244), .B(DATAIN[21]), .S(n154), .Z(n3135) );
  MUX2_X1 U1164 ( .A(n4243), .B(DATAIN[20]), .S(n154), .Z(n3134) );
  MUX2_X1 U1165 ( .A(n4242), .B(DATAIN[19]), .S(n154), .Z(n3133) );
  MUX2_X1 U1166 ( .A(n4241), .B(DATAIN[18]), .S(n154), .Z(n3132) );
  MUX2_X1 U1167 ( .A(n4240), .B(DATAIN[17]), .S(n154), .Z(n3131) );
  MUX2_X1 U1168 ( .A(n4239), .B(DATAIN[16]), .S(n154), .Z(n3130) );
  MUX2_X1 U1169 ( .A(n4238), .B(DATAIN[15]), .S(n154), .Z(n3129) );
  MUX2_X1 U1170 ( .A(n4237), .B(DATAIN[14]), .S(n154), .Z(n3128) );
  MUX2_X1 U1171 ( .A(n4236), .B(DATAIN[13]), .S(n154), .Z(n3127) );
  MUX2_X1 U1172 ( .A(n4235), .B(DATAIN[12]), .S(n154), .Z(n3126) );
  MUX2_X1 U1173 ( .A(n4234), .B(DATAIN[11]), .S(n153), .Z(n3125) );
  MUX2_X1 U1174 ( .A(n4233), .B(DATAIN[10]), .S(n153), .Z(n3124) );
  MUX2_X1 U1175 ( .A(n4232), .B(DATAIN[9]), .S(n153), .Z(n3123) );
  MUX2_X1 U1176 ( .A(n4231), .B(DATAIN[8]), .S(n153), .Z(n3122) );
  MUX2_X1 U1177 ( .A(n4230), .B(DATAIN[7]), .S(n153), .Z(n3121) );
  MUX2_X1 U1178 ( .A(n4229), .B(DATAIN[6]), .S(n153), .Z(n3120) );
  MUX2_X1 U1179 ( .A(n4228), .B(DATAIN[5]), .S(n153), .Z(n3119) );
  MUX2_X1 U1180 ( .A(n4227), .B(DATAIN[4]), .S(n153), .Z(n3118) );
  MUX2_X1 U1181 ( .A(n4226), .B(DATAIN[3]), .S(n153), .Z(n3117) );
  MUX2_X1 U1182 ( .A(n4225), .B(DATAIN[2]), .S(n153), .Z(n3116) );
  MUX2_X1 U1183 ( .A(n4224), .B(DATAIN[1]), .S(n153), .Z(n3115) );
  MUX2_X1 U1184 ( .A(n4223), .B(DATAIN[0]), .S(n153), .Z(n3114) );
  AND2_X1 U1185 ( .A1(n909), .A2(n870), .ZN(n1044) );
  MUX2_X1 U1186 ( .A(n4222), .B(DATAIN[31]), .S(n158), .Z(n3113) );
  MUX2_X1 U1187 ( .A(n4221), .B(DATAIN[30]), .S(n158), .Z(n3112) );
  MUX2_X1 U1188 ( .A(n4220), .B(DATAIN[29]), .S(n158), .Z(n3111) );
  MUX2_X1 U1189 ( .A(n4219), .B(DATAIN[28]), .S(n158), .Z(n3110) );
  MUX2_X1 U1190 ( .A(n4218), .B(DATAIN[27]), .S(n158), .Z(n3109) );
  MUX2_X1 U1191 ( .A(n4217), .B(DATAIN[26]), .S(n158), .Z(n3108) );
  MUX2_X1 U1192 ( .A(n4216), .B(DATAIN[25]), .S(n158), .Z(n3107) );
  MUX2_X1 U1193 ( .A(n4215), .B(DATAIN[24]), .S(n158), .Z(n3106) );
  MUX2_X1 U1194 ( .A(n4214), .B(DATAIN[23]), .S(n157), .Z(n3105) );
  MUX2_X1 U1195 ( .A(n4213), .B(DATAIN[22]), .S(n157), .Z(n3104) );
  MUX2_X1 U1196 ( .A(n4212), .B(DATAIN[21]), .S(n157), .Z(n3103) );
  MUX2_X1 U1197 ( .A(n4211), .B(DATAIN[20]), .S(n157), .Z(n3102) );
  MUX2_X1 U1198 ( .A(n4210), .B(DATAIN[19]), .S(n157), .Z(n3101) );
  MUX2_X1 U1199 ( .A(n4209), .B(DATAIN[18]), .S(n157), .Z(n3100) );
  MUX2_X1 U1200 ( .A(n4208), .B(DATAIN[17]), .S(n157), .Z(n3099) );
  MUX2_X1 U1201 ( .A(n4207), .B(DATAIN[16]), .S(n157), .Z(n3098) );
  MUX2_X1 U1202 ( .A(n4206), .B(DATAIN[15]), .S(n157), .Z(n3097) );
  MUX2_X1 U1203 ( .A(n4205), .B(DATAIN[14]), .S(n157), .Z(n3096) );
  MUX2_X1 U1204 ( .A(n4204), .B(DATAIN[13]), .S(n157), .Z(n3095) );
  MUX2_X1 U1205 ( .A(n4203), .B(DATAIN[12]), .S(n157), .Z(n3094) );
  MUX2_X1 U1206 ( .A(n4202), .B(DATAIN[11]), .S(n156), .Z(n3093) );
  MUX2_X1 U1207 ( .A(n4201), .B(DATAIN[10]), .S(n156), .Z(n3092) );
  MUX2_X1 U1208 ( .A(n4200), .B(DATAIN[9]), .S(n156), .Z(n3091) );
  MUX2_X1 U1209 ( .A(n4199), .B(DATAIN[8]), .S(n156), .Z(n3090) );
  MUX2_X1 U1210 ( .A(n4198), .B(DATAIN[7]), .S(n156), .Z(n3089) );
  MUX2_X1 U1211 ( .A(n4197), .B(DATAIN[6]), .S(n156), .Z(n3088) );
  MUX2_X1 U1212 ( .A(n4196), .B(DATAIN[5]), .S(n156), .Z(n3087) );
  MUX2_X1 U1213 ( .A(n4195), .B(DATAIN[4]), .S(n156), .Z(n3086) );
  MUX2_X1 U1214 ( .A(n4194), .B(DATAIN[3]), .S(n156), .Z(n3085) );
  MUX2_X1 U1215 ( .A(n4193), .B(DATAIN[2]), .S(n156), .Z(n3084) );
  MUX2_X1 U1216 ( .A(n4192), .B(DATAIN[1]), .S(n156), .Z(n3083) );
  MUX2_X1 U1217 ( .A(n4191), .B(DATAIN[0]), .S(n156), .Z(n3082) );
  AND2_X1 U1218 ( .A1(n909), .A2(n872), .ZN(n1045) );
  AND3_X1 U1219 ( .A1(n875), .A2(n874), .A3(ADD_WR[3]), .ZN(n909) );
  MUX2_X1 U1220 ( .A(n1046), .B(DATAIN[31]), .S(n161), .Z(n3081) );
  MUX2_X1 U1221 ( .A(n1048), .B(DATAIN[30]), .S(n161), .Z(n3080) );
  MUX2_X1 U1222 ( .A(n1049), .B(DATAIN[29]), .S(n161), .Z(n3079) );
  MUX2_X1 U1223 ( .A(n1050), .B(DATAIN[28]), .S(n161), .Z(n3078) );
  MUX2_X1 U1224 ( .A(n1051), .B(DATAIN[27]), .S(n161), .Z(n3077) );
  MUX2_X1 U1225 ( .A(n1052), .B(DATAIN[26]), .S(n161), .Z(n3076) );
  MUX2_X1 U1226 ( .A(n1053), .B(DATAIN[25]), .S(n161), .Z(n3075) );
  MUX2_X1 U1227 ( .A(n1054), .B(DATAIN[24]), .S(n161), .Z(n3074) );
  MUX2_X1 U1228 ( .A(n1055), .B(DATAIN[23]), .S(n160), .Z(n3073) );
  MUX2_X1 U1229 ( .A(n1056), .B(DATAIN[22]), .S(n160), .Z(n3072) );
  MUX2_X1 U1230 ( .A(n1057), .B(DATAIN[21]), .S(n160), .Z(n3071) );
  MUX2_X1 U1231 ( .A(n1058), .B(DATAIN[20]), .S(n160), .Z(n3070) );
  MUX2_X1 U1232 ( .A(n1059), .B(DATAIN[19]), .S(n160), .Z(n3069) );
  MUX2_X1 U1233 ( .A(n1060), .B(DATAIN[18]), .S(n160), .Z(n3068) );
  MUX2_X1 U1234 ( .A(n1061), .B(DATAIN[17]), .S(n160), .Z(n3067) );
  MUX2_X1 U1235 ( .A(n1062), .B(DATAIN[16]), .S(n160), .Z(n3066) );
  MUX2_X1 U1236 ( .A(n1063), .B(DATAIN[15]), .S(n160), .Z(n3065) );
  MUX2_X1 U1237 ( .A(n1064), .B(DATAIN[14]), .S(n160), .Z(n3064) );
  MUX2_X1 U1238 ( .A(n1065), .B(DATAIN[13]), .S(n160), .Z(n3063) );
  MUX2_X1 U1239 ( .A(n1066), .B(DATAIN[12]), .S(n160), .Z(n3062) );
  MUX2_X1 U1240 ( .A(n1067), .B(DATAIN[11]), .S(n159), .Z(n3061) );
  MUX2_X1 U1241 ( .A(n1068), .B(DATAIN[10]), .S(n159), .Z(n3060) );
  MUX2_X1 U1242 ( .A(n1069), .B(DATAIN[9]), .S(n159), .Z(n3059) );
  MUX2_X1 U1243 ( .A(n1070), .B(DATAIN[8]), .S(n159), .Z(n3058) );
  MUX2_X1 U1244 ( .A(n1071), .B(DATAIN[7]), .S(n159), .Z(n3057) );
  MUX2_X1 U1245 ( .A(n1072), .B(DATAIN[6]), .S(n159), .Z(n3056) );
  MUX2_X1 U1246 ( .A(n1073), .B(DATAIN[5]), .S(n159), .Z(n3055) );
  MUX2_X1 U1247 ( .A(n1074), .B(DATAIN[4]), .S(n159), .Z(n3054) );
  MUX2_X1 U1248 ( .A(n1075), .B(DATAIN[3]), .S(n159), .Z(n3053) );
  MUX2_X1 U1249 ( .A(n1076), .B(DATAIN[2]), .S(n159), .Z(n3052) );
  MUX2_X1 U1250 ( .A(n1077), .B(DATAIN[1]), .S(n159), .Z(n3051) );
  MUX2_X1 U1251 ( .A(n1078), .B(DATAIN[0]), .S(n159), .Z(n3050) );
  AND2_X1 U1252 ( .A1(n1079), .A2(n910), .ZN(n1047) );
  INV_X1 U1253 ( .A(n1080), .ZN(n3049) );
  MUX2_X1 U1254 ( .A(n517), .B(n593), .S(n164), .Z(n1080) );
  INV_X1 U1255 ( .A(n1082), .ZN(n3048) );
  MUX2_X1 U1256 ( .A(n518), .B(n592), .S(n164), .Z(n1082) );
  INV_X1 U1257 ( .A(n1083), .ZN(n3047) );
  MUX2_X1 U1258 ( .A(n519), .B(n591), .S(n164), .Z(n1083) );
  INV_X1 U1259 ( .A(n1084), .ZN(n3046) );
  MUX2_X1 U1260 ( .A(n520), .B(n590), .S(n164), .Z(n1084) );
  INV_X1 U1261 ( .A(n1085), .ZN(n3045) );
  MUX2_X1 U1262 ( .A(n521), .B(n589), .S(n164), .Z(n1085) );
  INV_X1 U1263 ( .A(n1086), .ZN(n3044) );
  MUX2_X1 U1264 ( .A(n522), .B(n588), .S(n164), .Z(n1086) );
  INV_X1 U1265 ( .A(n1087), .ZN(n3043) );
  MUX2_X1 U1266 ( .A(n523), .B(n587), .S(n164), .Z(n1087) );
  INV_X1 U1267 ( .A(n1088), .ZN(n3042) );
  MUX2_X1 U1268 ( .A(n524), .B(n586), .S(n164), .Z(n1088) );
  INV_X1 U1269 ( .A(n1089), .ZN(n3041) );
  MUX2_X1 U1270 ( .A(n525), .B(n585), .S(n163), .Z(n1089) );
  INV_X1 U1271 ( .A(n1090), .ZN(n3040) );
  MUX2_X1 U1272 ( .A(n526), .B(n584), .S(n163), .Z(n1090) );
  INV_X1 U1273 ( .A(n1091), .ZN(n3039) );
  MUX2_X1 U1274 ( .A(n527), .B(n583), .S(n163), .Z(n1091) );
  INV_X1 U1275 ( .A(n1092), .ZN(n3038) );
  MUX2_X1 U1276 ( .A(n528), .B(n582), .S(n163), .Z(n1092) );
  INV_X1 U1277 ( .A(n1093), .ZN(n3037) );
  MUX2_X1 U1278 ( .A(n529), .B(n581), .S(n163), .Z(n1093) );
  INV_X1 U1279 ( .A(n1094), .ZN(n3036) );
  MUX2_X1 U1280 ( .A(n530), .B(n580), .S(n163), .Z(n1094) );
  INV_X1 U1281 ( .A(n1095), .ZN(n3035) );
  MUX2_X1 U1282 ( .A(n531), .B(n579), .S(n163), .Z(n1095) );
  INV_X1 U1283 ( .A(n1096), .ZN(n3034) );
  MUX2_X1 U1284 ( .A(n532), .B(n578), .S(n163), .Z(n1096) );
  INV_X1 U1285 ( .A(n1097), .ZN(n3033) );
  MUX2_X1 U1286 ( .A(n533), .B(n577), .S(n163), .Z(n1097) );
  INV_X1 U1287 ( .A(n1098), .ZN(n3032) );
  MUX2_X1 U1288 ( .A(n534), .B(n576), .S(n163), .Z(n1098) );
  INV_X1 U1289 ( .A(n1099), .ZN(n3031) );
  MUX2_X1 U1290 ( .A(n535), .B(n575), .S(n163), .Z(n1099) );
  INV_X1 U1291 ( .A(n1100), .ZN(n3030) );
  MUX2_X1 U1292 ( .A(n536), .B(n574), .S(n163), .Z(n1100) );
  INV_X1 U1293 ( .A(n1101), .ZN(n3029) );
  MUX2_X1 U1294 ( .A(n537), .B(n573), .S(n162), .Z(n1101) );
  INV_X1 U1295 ( .A(n1102), .ZN(n3028) );
  MUX2_X1 U1296 ( .A(n538), .B(n572), .S(n162), .Z(n1102) );
  INV_X1 U1297 ( .A(n1103), .ZN(n3027) );
  MUX2_X1 U1298 ( .A(n539), .B(n571), .S(n162), .Z(n1103) );
  INV_X1 U1299 ( .A(n1104), .ZN(n3026) );
  MUX2_X1 U1300 ( .A(n540), .B(n570), .S(n162), .Z(n1104) );
  INV_X1 U1301 ( .A(n1105), .ZN(n3025) );
  MUX2_X1 U1302 ( .A(n541), .B(n569), .S(n162), .Z(n1105) );
  INV_X1 U1303 ( .A(n1106), .ZN(n3024) );
  MUX2_X1 U1304 ( .A(n542), .B(n568), .S(n162), .Z(n1106) );
  INV_X1 U1305 ( .A(n1107), .ZN(n3023) );
  MUX2_X1 U1306 ( .A(n543), .B(n567), .S(n162), .Z(n1107) );
  INV_X1 U1307 ( .A(n1108), .ZN(n3022) );
  MUX2_X1 U1308 ( .A(n544), .B(n566), .S(n162), .Z(n1108) );
  INV_X1 U1309 ( .A(n1109), .ZN(n3021) );
  MUX2_X1 U1310 ( .A(n545), .B(n565), .S(n162), .Z(n1109) );
  INV_X1 U1311 ( .A(n1110), .ZN(n3020) );
  MUX2_X1 U1312 ( .A(n546), .B(n564), .S(n162), .Z(n1110) );
  INV_X1 U1313 ( .A(n1111), .ZN(n3019) );
  MUX2_X1 U1314 ( .A(n547), .B(n563), .S(n162), .Z(n1111) );
  INV_X1 U1315 ( .A(n1112), .ZN(n3018) );
  MUX2_X1 U1316 ( .A(n548), .B(n562), .S(n162), .Z(n1112) );
  AND2_X1 U1317 ( .A1(n1079), .A2(n763), .ZN(n1081) );
  MUX2_X1 U1318 ( .A(n4190), .B(DATAIN[31]), .S(n167), .Z(n3017) );
  MUX2_X1 U1319 ( .A(n4189), .B(DATAIN[30]), .S(n167), .Z(n3016) );
  MUX2_X1 U1320 ( .A(n4188), .B(DATAIN[29]), .S(n167), .Z(n3015) );
  MUX2_X1 U1321 ( .A(n4187), .B(DATAIN[28]), .S(n167), .Z(n3014) );
  MUX2_X1 U1322 ( .A(n4186), .B(DATAIN[27]), .S(n167), .Z(n3013) );
  MUX2_X1 U1323 ( .A(n4185), .B(DATAIN[26]), .S(n167), .Z(n3012) );
  MUX2_X1 U1324 ( .A(n4184), .B(DATAIN[25]), .S(n167), .Z(n3011) );
  MUX2_X1 U1325 ( .A(n4183), .B(DATAIN[24]), .S(n167), .Z(n3010) );
  MUX2_X1 U1326 ( .A(n4182), .B(DATAIN[23]), .S(n166), .Z(n3009) );
  MUX2_X1 U1327 ( .A(n4181), .B(DATAIN[22]), .S(n166), .Z(n3008) );
  MUX2_X1 U1328 ( .A(n4180), .B(DATAIN[21]), .S(n166), .Z(n3007) );
  MUX2_X1 U1329 ( .A(n4179), .B(DATAIN[20]), .S(n166), .Z(n3006) );
  MUX2_X1 U1330 ( .A(n4178), .B(DATAIN[19]), .S(n166), .Z(n3005) );
  MUX2_X1 U1331 ( .A(n4177), .B(DATAIN[18]), .S(n166), .Z(n3004) );
  MUX2_X1 U1332 ( .A(n4176), .B(DATAIN[17]), .S(n166), .Z(n3003) );
  MUX2_X1 U1333 ( .A(n4175), .B(DATAIN[16]), .S(n166), .Z(n3002) );
  MUX2_X1 U1334 ( .A(n4174), .B(DATAIN[15]), .S(n166), .Z(n3001) );
  MUX2_X1 U1335 ( .A(n4173), .B(DATAIN[14]), .S(n166), .Z(n3000) );
  MUX2_X1 U1336 ( .A(n4172), .B(DATAIN[13]), .S(n166), .Z(n2999) );
  MUX2_X1 U1337 ( .A(n4171), .B(DATAIN[12]), .S(n166), .Z(n2998) );
  MUX2_X1 U1338 ( .A(n4170), .B(DATAIN[11]), .S(n165), .Z(n2997) );
  MUX2_X1 U1339 ( .A(n4169), .B(DATAIN[10]), .S(n165), .Z(n2996) );
  MUX2_X1 U1340 ( .A(n4168), .B(DATAIN[9]), .S(n165), .Z(n2995) );
  MUX2_X1 U1341 ( .A(n4167), .B(DATAIN[8]), .S(n165), .Z(n2994) );
  MUX2_X1 U1342 ( .A(n4166), .B(DATAIN[7]), .S(n165), .Z(n2993) );
  MUX2_X1 U1343 ( .A(n4165), .B(DATAIN[6]), .S(n165), .Z(n2992) );
  MUX2_X1 U1344 ( .A(n4164), .B(DATAIN[5]), .S(n165), .Z(n2991) );
  MUX2_X1 U1345 ( .A(n4163), .B(DATAIN[4]), .S(n165), .Z(n2990) );
  MUX2_X1 U1346 ( .A(n4162), .B(DATAIN[3]), .S(n165), .Z(n2989) );
  MUX2_X1 U1347 ( .A(n4161), .B(DATAIN[2]), .S(n165), .Z(n2988) );
  MUX2_X1 U1348 ( .A(n4160), .B(DATAIN[1]), .S(n165), .Z(n2987) );
  MUX2_X1 U1349 ( .A(n4159), .B(DATAIN[0]), .S(n165), .Z(n2986) );
  AND2_X1 U1350 ( .A1(n1079), .A2(n766), .ZN(n1113) );
  MUX2_X1 U1351 ( .A(n4158), .B(DATAIN[31]), .S(n170), .Z(n2985) );
  MUX2_X1 U1352 ( .A(n4157), .B(DATAIN[30]), .S(n170), .Z(n2984) );
  MUX2_X1 U1353 ( .A(n4156), .B(DATAIN[29]), .S(n170), .Z(n2983) );
  MUX2_X1 U1354 ( .A(n4155), .B(DATAIN[28]), .S(n170), .Z(n2982) );
  MUX2_X1 U1355 ( .A(n4154), .B(DATAIN[27]), .S(n170), .Z(n2981) );
  MUX2_X1 U1356 ( .A(n4153), .B(DATAIN[26]), .S(n170), .Z(n2980) );
  MUX2_X1 U1357 ( .A(n4152), .B(DATAIN[25]), .S(n170), .Z(n2979) );
  MUX2_X1 U1358 ( .A(n4151), .B(DATAIN[24]), .S(n170), .Z(n2978) );
  MUX2_X1 U1359 ( .A(n4150), .B(DATAIN[23]), .S(n169), .Z(n2977) );
  MUX2_X1 U1360 ( .A(n4149), .B(DATAIN[22]), .S(n169), .Z(n2976) );
  MUX2_X1 U1361 ( .A(n4148), .B(DATAIN[21]), .S(n169), .Z(n2975) );
  MUX2_X1 U1362 ( .A(n4147), .B(DATAIN[20]), .S(n169), .Z(n2974) );
  MUX2_X1 U1363 ( .A(n4146), .B(DATAIN[19]), .S(n169), .Z(n2973) );
  MUX2_X1 U1364 ( .A(n4145), .B(DATAIN[18]), .S(n169), .Z(n2972) );
  MUX2_X1 U1365 ( .A(n4144), .B(DATAIN[17]), .S(n169), .Z(n2971) );
  MUX2_X1 U1366 ( .A(n4143), .B(DATAIN[16]), .S(n169), .Z(n2970) );
  MUX2_X1 U1367 ( .A(n4142), .B(DATAIN[15]), .S(n169), .Z(n2969) );
  MUX2_X1 U1368 ( .A(n4141), .B(DATAIN[14]), .S(n169), .Z(n2968) );
  MUX2_X1 U1369 ( .A(n4140), .B(DATAIN[13]), .S(n169), .Z(n2967) );
  MUX2_X1 U1370 ( .A(n4139), .B(DATAIN[12]), .S(n169), .Z(n2966) );
  MUX2_X1 U1371 ( .A(n4138), .B(DATAIN[11]), .S(n168), .Z(n2965) );
  MUX2_X1 U1372 ( .A(n4137), .B(DATAIN[10]), .S(n168), .Z(n2964) );
  MUX2_X1 U1373 ( .A(n4136), .B(DATAIN[9]), .S(n168), .Z(n2963) );
  MUX2_X1 U1374 ( .A(n4135), .B(DATAIN[8]), .S(n168), .Z(n2962) );
  MUX2_X1 U1375 ( .A(n4134), .B(DATAIN[7]), .S(n168), .Z(n2961) );
  MUX2_X1 U1376 ( .A(n4133), .B(DATAIN[6]), .S(n168), .Z(n2960) );
  MUX2_X1 U1377 ( .A(n4132), .B(DATAIN[5]), .S(n168), .Z(n2959) );
  MUX2_X1 U1378 ( .A(n4131), .B(DATAIN[4]), .S(n168), .Z(n2958) );
  MUX2_X1 U1379 ( .A(n4130), .B(DATAIN[3]), .S(n168), .Z(n2957) );
  MUX2_X1 U1380 ( .A(n4129), .B(DATAIN[2]), .S(n168), .Z(n2956) );
  MUX2_X1 U1381 ( .A(n4128), .B(DATAIN[1]), .S(n168), .Z(n2955) );
  MUX2_X1 U1382 ( .A(n4127), .B(DATAIN[0]), .S(n168), .Z(n2954) );
  AND2_X1 U1383 ( .A1(n1079), .A2(n768), .ZN(n1114) );
  INV_X1 U1384 ( .A(n1115), .ZN(n2953) );
  MUX2_X1 U1385 ( .A(n613), .B(n593), .S(n173), .Z(n1115) );
  INV_X1 U1386 ( .A(n1117), .ZN(n2952) );
  MUX2_X1 U1387 ( .A(n614), .B(n592), .S(n173), .Z(n1117) );
  INV_X1 U1388 ( .A(n1118), .ZN(n2951) );
  MUX2_X1 U1389 ( .A(n615), .B(n591), .S(n173), .Z(n1118) );
  INV_X1 U1390 ( .A(n1119), .ZN(n2950) );
  MUX2_X1 U1391 ( .A(n616), .B(n590), .S(n173), .Z(n1119) );
  INV_X1 U1392 ( .A(n1120), .ZN(n2949) );
  MUX2_X1 U1393 ( .A(n617), .B(n589), .S(n173), .Z(n1120) );
  INV_X1 U1394 ( .A(n1121), .ZN(n2948) );
  MUX2_X1 U1395 ( .A(n618), .B(n588), .S(n173), .Z(n1121) );
  INV_X1 U1396 ( .A(n1122), .ZN(n2947) );
  MUX2_X1 U1397 ( .A(n619), .B(n587), .S(n173), .Z(n1122) );
  INV_X1 U1398 ( .A(n1123), .ZN(n2946) );
  MUX2_X1 U1399 ( .A(n620), .B(n586), .S(n173), .Z(n1123) );
  INV_X1 U1400 ( .A(n1124), .ZN(n2945) );
  MUX2_X1 U1401 ( .A(n621), .B(n585), .S(n172), .Z(n1124) );
  INV_X1 U1402 ( .A(n1125), .ZN(n2944) );
  MUX2_X1 U1403 ( .A(n622), .B(n584), .S(n172), .Z(n1125) );
  INV_X1 U1404 ( .A(n1126), .ZN(n2943) );
  MUX2_X1 U1405 ( .A(n623), .B(n583), .S(n172), .Z(n1126) );
  INV_X1 U1406 ( .A(n1127), .ZN(n2942) );
  MUX2_X1 U1407 ( .A(n624), .B(n582), .S(n172), .Z(n1127) );
  INV_X1 U1408 ( .A(n1128), .ZN(n2941) );
  MUX2_X1 U1409 ( .A(n625), .B(n581), .S(n172), .Z(n1128) );
  INV_X1 U1410 ( .A(n1129), .ZN(n2940) );
  MUX2_X1 U1411 ( .A(n626), .B(n580), .S(n172), .Z(n1129) );
  INV_X1 U1412 ( .A(n1130), .ZN(n2939) );
  MUX2_X1 U1413 ( .A(n627), .B(n579), .S(n172), .Z(n1130) );
  INV_X1 U1414 ( .A(n1131), .ZN(n2938) );
  MUX2_X1 U1415 ( .A(n628), .B(n578), .S(n172), .Z(n1131) );
  INV_X1 U1416 ( .A(n1132), .ZN(n2937) );
  MUX2_X1 U1417 ( .A(n629), .B(n577), .S(n172), .Z(n1132) );
  INV_X1 U1418 ( .A(n1133), .ZN(n2936) );
  MUX2_X1 U1419 ( .A(n630), .B(n576), .S(n172), .Z(n1133) );
  INV_X1 U1420 ( .A(n1134), .ZN(n2935) );
  MUX2_X1 U1421 ( .A(n631), .B(n575), .S(n172), .Z(n1134) );
  INV_X1 U1422 ( .A(n1135), .ZN(n2934) );
  MUX2_X1 U1423 ( .A(n632), .B(n574), .S(n172), .Z(n1135) );
  INV_X1 U1424 ( .A(n1136), .ZN(n2933) );
  MUX2_X1 U1425 ( .A(n633), .B(n573), .S(n171), .Z(n1136) );
  INV_X1 U1426 ( .A(n1137), .ZN(n2932) );
  MUX2_X1 U1427 ( .A(n634), .B(n572), .S(n171), .Z(n1137) );
  INV_X1 U1428 ( .A(n1138), .ZN(n2931) );
  MUX2_X1 U1429 ( .A(n635), .B(n571), .S(n171), .Z(n1138) );
  INV_X1 U1430 ( .A(n1139), .ZN(n2930) );
  MUX2_X1 U1431 ( .A(n636), .B(n570), .S(n171), .Z(n1139) );
  INV_X1 U1432 ( .A(n1140), .ZN(n2929) );
  MUX2_X1 U1433 ( .A(n637), .B(n569), .S(n171), .Z(n1140) );
  INV_X1 U1434 ( .A(n1141), .ZN(n2928) );
  MUX2_X1 U1435 ( .A(n638), .B(n568), .S(n171), .Z(n1141) );
  INV_X1 U1436 ( .A(n1142), .ZN(n2927) );
  MUX2_X1 U1437 ( .A(n639), .B(n567), .S(n171), .Z(n1142) );
  INV_X1 U1438 ( .A(n1143), .ZN(n2926) );
  MUX2_X1 U1439 ( .A(n640), .B(n566), .S(n171), .Z(n1143) );
  INV_X1 U1440 ( .A(n1144), .ZN(n2925) );
  MUX2_X1 U1441 ( .A(n641), .B(n565), .S(n171), .Z(n1144) );
  INV_X1 U1442 ( .A(n1145), .ZN(n2924) );
  MUX2_X1 U1443 ( .A(n642), .B(n564), .S(n171), .Z(n1145) );
  INV_X1 U1444 ( .A(n1146), .ZN(n2923) );
  MUX2_X1 U1445 ( .A(n643), .B(n563), .S(n171), .Z(n1146) );
  INV_X1 U1446 ( .A(n1147), .ZN(n2922) );
  MUX2_X1 U1447 ( .A(n644), .B(n562), .S(n171), .Z(n1147) );
  AND2_X1 U1448 ( .A1(n1079), .A2(n802), .ZN(n1116) );
  MUX2_X1 U1449 ( .A(n1148), .B(DATAIN[31]), .S(n176), .Z(n2921) );
  MUX2_X1 U1450 ( .A(n1150), .B(DATAIN[30]), .S(n176), .Z(n2920) );
  MUX2_X1 U1451 ( .A(n1151), .B(DATAIN[29]), .S(n176), .Z(n2919) );
  MUX2_X1 U1452 ( .A(n1152), .B(DATAIN[28]), .S(n176), .Z(n2918) );
  MUX2_X1 U1453 ( .A(n1153), .B(DATAIN[27]), .S(n176), .Z(n2917) );
  MUX2_X1 U1454 ( .A(n1154), .B(DATAIN[26]), .S(n176), .Z(n2916) );
  MUX2_X1 U1455 ( .A(n1155), .B(DATAIN[25]), .S(n176), .Z(n2915) );
  MUX2_X1 U1456 ( .A(n1156), .B(DATAIN[24]), .S(n176), .Z(n2914) );
  MUX2_X1 U1457 ( .A(n1157), .B(DATAIN[23]), .S(n175), .Z(n2913) );
  MUX2_X1 U1458 ( .A(n1158), .B(DATAIN[22]), .S(n175), .Z(n2912) );
  MUX2_X1 U1459 ( .A(n1159), .B(DATAIN[21]), .S(n175), .Z(n2911) );
  MUX2_X1 U1460 ( .A(n1160), .B(DATAIN[20]), .S(n175), .Z(n2910) );
  MUX2_X1 U1461 ( .A(n1161), .B(DATAIN[19]), .S(n175), .Z(n2909) );
  MUX2_X1 U1462 ( .A(n1162), .B(DATAIN[18]), .S(n175), .Z(n2908) );
  MUX2_X1 U1463 ( .A(n1163), .B(DATAIN[17]), .S(n175), .Z(n2907) );
  MUX2_X1 U1464 ( .A(n1164), .B(DATAIN[16]), .S(n175), .Z(n2906) );
  MUX2_X1 U1465 ( .A(n1165), .B(DATAIN[15]), .S(n175), .Z(n2905) );
  MUX2_X1 U1466 ( .A(n1166), .B(DATAIN[14]), .S(n175), .Z(n2904) );
  MUX2_X1 U1467 ( .A(n1167), .B(DATAIN[13]), .S(n175), .Z(n2903) );
  MUX2_X1 U1468 ( .A(n1168), .B(DATAIN[12]), .S(n175), .Z(n2902) );
  MUX2_X1 U1469 ( .A(n1169), .B(DATAIN[11]), .S(n174), .Z(n2901) );
  MUX2_X1 U1470 ( .A(n1170), .B(DATAIN[10]), .S(n174), .Z(n2900) );
  MUX2_X1 U1471 ( .A(n1171), .B(DATAIN[9]), .S(n174), .Z(n2899) );
  MUX2_X1 U1472 ( .A(n1172), .B(DATAIN[8]), .S(n174), .Z(n2898) );
  MUX2_X1 U1473 ( .A(n1173), .B(DATAIN[7]), .S(n174), .Z(n2897) );
  MUX2_X1 U1474 ( .A(n1174), .B(DATAIN[6]), .S(n174), .Z(n2896) );
  MUX2_X1 U1475 ( .A(n1175), .B(DATAIN[5]), .S(n174), .Z(n2895) );
  MUX2_X1 U1476 ( .A(n1176), .B(DATAIN[4]), .S(n174), .Z(n2894) );
  MUX2_X1 U1477 ( .A(n1177), .B(DATAIN[3]), .S(n174), .Z(n2893) );
  MUX2_X1 U1478 ( .A(n1178), .B(DATAIN[2]), .S(n174), .Z(n2892) );
  MUX2_X1 U1479 ( .A(n1179), .B(DATAIN[1]), .S(n174), .Z(n2891) );
  MUX2_X1 U1480 ( .A(n1180), .B(DATAIN[0]), .S(n174), .Z(n2890) );
  AND2_X1 U1481 ( .A1(n1079), .A2(n836), .ZN(n1149) );
  MUX2_X1 U1482 ( .A(n4126), .B(DATAIN[31]), .S(n179), .Z(n2889) );
  MUX2_X1 U1483 ( .A(n4125), .B(DATAIN[30]), .S(n179), .Z(n2888) );
  MUX2_X1 U1484 ( .A(n4124), .B(DATAIN[29]), .S(n179), .Z(n2887) );
  MUX2_X1 U1485 ( .A(n4123), .B(DATAIN[28]), .S(n179), .Z(n2886) );
  MUX2_X1 U1486 ( .A(n4122), .B(DATAIN[27]), .S(n179), .Z(n2885) );
  MUX2_X1 U1487 ( .A(n4121), .B(DATAIN[26]), .S(n179), .Z(n2884) );
  MUX2_X1 U1488 ( .A(n4120), .B(DATAIN[25]), .S(n179), .Z(n2883) );
  MUX2_X1 U1489 ( .A(n4119), .B(DATAIN[24]), .S(n179), .Z(n2882) );
  MUX2_X1 U1490 ( .A(n4118), .B(DATAIN[23]), .S(n178), .Z(n2881) );
  MUX2_X1 U1491 ( .A(n4117), .B(DATAIN[22]), .S(n178), .Z(n2880) );
  MUX2_X1 U1492 ( .A(n4116), .B(DATAIN[21]), .S(n178), .Z(n2879) );
  MUX2_X1 U1493 ( .A(n4115), .B(DATAIN[20]), .S(n178), .Z(n2878) );
  MUX2_X1 U1494 ( .A(n4114), .B(DATAIN[19]), .S(n178), .Z(n2877) );
  MUX2_X1 U1495 ( .A(n4113), .B(DATAIN[18]), .S(n178), .Z(n2876) );
  MUX2_X1 U1496 ( .A(n4112), .B(DATAIN[17]), .S(n178), .Z(n2875) );
  MUX2_X1 U1497 ( .A(n4111), .B(DATAIN[16]), .S(n178), .Z(n2874) );
  MUX2_X1 U1498 ( .A(n4110), .B(DATAIN[15]), .S(n178), .Z(n2873) );
  MUX2_X1 U1499 ( .A(n4109), .B(DATAIN[14]), .S(n178), .Z(n2872) );
  MUX2_X1 U1500 ( .A(n4108), .B(DATAIN[13]), .S(n178), .Z(n2871) );
  MUX2_X1 U1501 ( .A(n4107), .B(DATAIN[12]), .S(n178), .Z(n2870) );
  MUX2_X1 U1502 ( .A(n4106), .B(DATAIN[11]), .S(n177), .Z(n2869) );
  MUX2_X1 U1503 ( .A(n4105), .B(DATAIN[10]), .S(n177), .Z(n2868) );
  MUX2_X1 U1504 ( .A(n4104), .B(DATAIN[9]), .S(n177), .Z(n2867) );
  MUX2_X1 U1505 ( .A(n4103), .B(DATAIN[8]), .S(n177), .Z(n2866) );
  MUX2_X1 U1506 ( .A(n4102), .B(DATAIN[7]), .S(n177), .Z(n2865) );
  MUX2_X1 U1507 ( .A(n4101), .B(DATAIN[6]), .S(n177), .Z(n2864) );
  MUX2_X1 U1508 ( .A(n4100), .B(DATAIN[5]), .S(n177), .Z(n2863) );
  MUX2_X1 U1509 ( .A(n4099), .B(DATAIN[4]), .S(n177), .Z(n2862) );
  MUX2_X1 U1510 ( .A(n4098), .B(DATAIN[3]), .S(n177), .Z(n2861) );
  MUX2_X1 U1511 ( .A(n4097), .B(DATAIN[2]), .S(n177), .Z(n2860) );
  MUX2_X1 U1512 ( .A(n4096), .B(DATAIN[1]), .S(n177), .Z(n2859) );
  MUX2_X1 U1513 ( .A(n4095), .B(DATAIN[0]), .S(n177), .Z(n2858) );
  AND2_X1 U1514 ( .A1(n1079), .A2(n870), .ZN(n1181) );
  MUX2_X1 U1515 ( .A(n4094), .B(DATAIN[31]), .S(n182), .Z(n2857) );
  MUX2_X1 U1516 ( .A(n4093), .B(DATAIN[30]), .S(n182), .Z(n2856) );
  MUX2_X1 U1517 ( .A(n4092), .B(DATAIN[29]), .S(n182), .Z(n2855) );
  MUX2_X1 U1518 ( .A(n4091), .B(DATAIN[28]), .S(n182), .Z(n2854) );
  MUX2_X1 U1519 ( .A(n4090), .B(DATAIN[27]), .S(n182), .Z(n2853) );
  MUX2_X1 U1520 ( .A(n4089), .B(DATAIN[26]), .S(n182), .Z(n2852) );
  MUX2_X1 U1521 ( .A(n4088), .B(DATAIN[25]), .S(n182), .Z(n2851) );
  MUX2_X1 U1522 ( .A(n4087), .B(DATAIN[24]), .S(n182), .Z(n2850) );
  MUX2_X1 U1523 ( .A(n4086), .B(DATAIN[23]), .S(n181), .Z(n2849) );
  MUX2_X1 U1524 ( .A(n4085), .B(DATAIN[22]), .S(n181), .Z(n2848) );
  MUX2_X1 U1525 ( .A(n4084), .B(DATAIN[21]), .S(n181), .Z(n2847) );
  MUX2_X1 U1526 ( .A(n4083), .B(DATAIN[20]), .S(n181), .Z(n2846) );
  MUX2_X1 U1527 ( .A(n4082), .B(DATAIN[19]), .S(n181), .Z(n2845) );
  MUX2_X1 U1528 ( .A(n4081), .B(DATAIN[18]), .S(n181), .Z(n2844) );
  MUX2_X1 U1529 ( .A(n4080), .B(DATAIN[17]), .S(n181), .Z(n2843) );
  MUX2_X1 U1530 ( .A(n4079), .B(DATAIN[16]), .S(n181), .Z(n2842) );
  MUX2_X1 U1531 ( .A(n4078), .B(DATAIN[15]), .S(n181), .Z(n2841) );
  MUX2_X1 U1532 ( .A(n4077), .B(DATAIN[14]), .S(n181), .Z(n2840) );
  MUX2_X1 U1533 ( .A(n4076), .B(DATAIN[13]), .S(n181), .Z(n2839) );
  MUX2_X1 U1534 ( .A(n4075), .B(DATAIN[12]), .S(n181), .Z(n2838) );
  MUX2_X1 U1535 ( .A(n4074), .B(DATAIN[11]), .S(n180), .Z(n2837) );
  MUX2_X1 U1536 ( .A(n4073), .B(DATAIN[10]), .S(n180), .Z(n2836) );
  MUX2_X1 U1537 ( .A(n4072), .B(DATAIN[9]), .S(n180), .Z(n2835) );
  MUX2_X1 U1538 ( .A(n4071), .B(DATAIN[8]), .S(n180), .Z(n2834) );
  MUX2_X1 U1539 ( .A(n4070), .B(DATAIN[7]), .S(n180), .Z(n2833) );
  MUX2_X1 U1540 ( .A(n4069), .B(DATAIN[6]), .S(n180), .Z(n2832) );
  MUX2_X1 U1541 ( .A(n4068), .B(DATAIN[5]), .S(n180), .Z(n2831) );
  MUX2_X1 U1542 ( .A(n4067), .B(DATAIN[4]), .S(n180), .Z(n2830) );
  MUX2_X1 U1543 ( .A(n4066), .B(DATAIN[3]), .S(n180), .Z(n2829) );
  MUX2_X1 U1544 ( .A(n4065), .B(DATAIN[2]), .S(n180), .Z(n2828) );
  MUX2_X1 U1545 ( .A(n4064), .B(DATAIN[1]), .S(n180), .Z(n2827) );
  MUX2_X1 U1546 ( .A(n4063), .B(DATAIN[0]), .S(n180), .Z(n2826) );
  AND2_X1 U1547 ( .A1(n1079), .A2(n872), .ZN(n1182) );
  AND3_X1 U1548 ( .A1(n875), .A2(n873), .A3(ADD_WR[4]), .ZN(n1079) );
  MUX2_X1 U1549 ( .A(n4062), .B(DATAIN[31]), .S(n185), .Z(n2825) );
  MUX2_X1 U1550 ( .A(n4061), .B(DATAIN[30]), .S(n185), .Z(n2824) );
  MUX2_X1 U1551 ( .A(n4060), .B(DATAIN[29]), .S(n185), .Z(n2823) );
  MUX2_X1 U1552 ( .A(n4059), .B(DATAIN[28]), .S(n185), .Z(n2822) );
  MUX2_X1 U1553 ( .A(n4058), .B(DATAIN[27]), .S(n185), .Z(n2821) );
  MUX2_X1 U1554 ( .A(n4057), .B(DATAIN[26]), .S(n185), .Z(n2820) );
  MUX2_X1 U1555 ( .A(n4056), .B(DATAIN[25]), .S(n185), .Z(n2819) );
  MUX2_X1 U1556 ( .A(n4055), .B(DATAIN[24]), .S(n185), .Z(n2818) );
  MUX2_X1 U1557 ( .A(n4054), .B(DATAIN[23]), .S(n184), .Z(n2817) );
  MUX2_X1 U1558 ( .A(n4053), .B(DATAIN[22]), .S(n184), .Z(n2816) );
  MUX2_X1 U1559 ( .A(n4052), .B(DATAIN[21]), .S(n184), .Z(n2815) );
  MUX2_X1 U1560 ( .A(n4051), .B(DATAIN[20]), .S(n184), .Z(n2814) );
  MUX2_X1 U1561 ( .A(n4050), .B(DATAIN[19]), .S(n184), .Z(n2813) );
  MUX2_X1 U1562 ( .A(n4049), .B(DATAIN[18]), .S(n184), .Z(n2812) );
  MUX2_X1 U1563 ( .A(n4048), .B(DATAIN[17]), .S(n184), .Z(n2811) );
  MUX2_X1 U1564 ( .A(n4047), .B(DATAIN[16]), .S(n184), .Z(n2810) );
  MUX2_X1 U1565 ( .A(n4046), .B(DATAIN[15]), .S(n184), .Z(n2809) );
  MUX2_X1 U1566 ( .A(n4045), .B(DATAIN[14]), .S(n184), .Z(n2808) );
  MUX2_X1 U1567 ( .A(n4044), .B(DATAIN[13]), .S(n184), .Z(n2807) );
  MUX2_X1 U1568 ( .A(n4043), .B(DATAIN[12]), .S(n184), .Z(n2806) );
  MUX2_X1 U1569 ( .A(n4042), .B(DATAIN[11]), .S(n183), .Z(n2805) );
  MUX2_X1 U1570 ( .A(n4041), .B(DATAIN[10]), .S(n183), .Z(n2804) );
  MUX2_X1 U1571 ( .A(n4040), .B(DATAIN[9]), .S(n183), .Z(n2803) );
  MUX2_X1 U1572 ( .A(n4039), .B(DATAIN[8]), .S(n183), .Z(n2802) );
  MUX2_X1 U1573 ( .A(n4038), .B(DATAIN[7]), .S(n183), .Z(n2801) );
  MUX2_X1 U1574 ( .A(n4037), .B(DATAIN[6]), .S(n183), .Z(n2800) );
  MUX2_X1 U1575 ( .A(n4036), .B(DATAIN[5]), .S(n183), .Z(n2799) );
  MUX2_X1 U1576 ( .A(n4035), .B(DATAIN[4]), .S(n183), .Z(n2798) );
  MUX2_X1 U1577 ( .A(n4034), .B(DATAIN[3]), .S(n183), .Z(n2797) );
  MUX2_X1 U1578 ( .A(n4033), .B(DATAIN[2]), .S(n183), .Z(n2796) );
  MUX2_X1 U1579 ( .A(n4032), .B(DATAIN[1]), .S(n183), .Z(n2795) );
  MUX2_X1 U1580 ( .A(n4031), .B(DATAIN[0]), .S(n183), .Z(n2794) );
  AND2_X1 U1581 ( .A1(n1184), .A2(n910), .ZN(n1183) );
  MUX2_X1 U1582 ( .A(n4030), .B(DATAIN[31]), .S(n188), .Z(n2793) );
  MUX2_X1 U1583 ( .A(n4029), .B(DATAIN[30]), .S(n188), .Z(n2792) );
  MUX2_X1 U1584 ( .A(n4028), .B(DATAIN[29]), .S(n188), .Z(n2791) );
  MUX2_X1 U1585 ( .A(n4027), .B(DATAIN[28]), .S(n188), .Z(n2790) );
  MUX2_X1 U1586 ( .A(n4026), .B(DATAIN[27]), .S(n188), .Z(n2789) );
  MUX2_X1 U1587 ( .A(n4025), .B(DATAIN[26]), .S(n188), .Z(n2788) );
  MUX2_X1 U1588 ( .A(n4024), .B(DATAIN[25]), .S(n188), .Z(n2787) );
  MUX2_X1 U1589 ( .A(n4023), .B(DATAIN[24]), .S(n188), .Z(n2786) );
  MUX2_X1 U1590 ( .A(n4022), .B(DATAIN[23]), .S(n187), .Z(n2785) );
  MUX2_X1 U1591 ( .A(n4021), .B(DATAIN[22]), .S(n187), .Z(n2784) );
  MUX2_X1 U1592 ( .A(n4020), .B(DATAIN[21]), .S(n187), .Z(n2783) );
  MUX2_X1 U1593 ( .A(n4019), .B(DATAIN[20]), .S(n187), .Z(n2782) );
  MUX2_X1 U1594 ( .A(n4018), .B(DATAIN[19]), .S(n187), .Z(n2781) );
  MUX2_X1 U1595 ( .A(n4017), .B(DATAIN[18]), .S(n187), .Z(n2780) );
  MUX2_X1 U1596 ( .A(n4016), .B(DATAIN[17]), .S(n187), .Z(n2779) );
  MUX2_X1 U1597 ( .A(n4015), .B(DATAIN[16]), .S(n187), .Z(n2778) );
  MUX2_X1 U1598 ( .A(n4014), .B(DATAIN[15]), .S(n187), .Z(n2777) );
  MUX2_X1 U1599 ( .A(n4013), .B(DATAIN[14]), .S(n187), .Z(n2776) );
  MUX2_X1 U1600 ( .A(n4012), .B(DATAIN[13]), .S(n187), .Z(n2775) );
  MUX2_X1 U1601 ( .A(n4011), .B(DATAIN[12]), .S(n187), .Z(n2774) );
  MUX2_X1 U1602 ( .A(n4010), .B(DATAIN[11]), .S(n186), .Z(n2773) );
  MUX2_X1 U1603 ( .A(n4009), .B(DATAIN[10]), .S(n186), .Z(n2772) );
  MUX2_X1 U1604 ( .A(n4008), .B(DATAIN[9]), .S(n186), .Z(n2771) );
  MUX2_X1 U1605 ( .A(n4007), .B(DATAIN[8]), .S(n186), .Z(n2770) );
  MUX2_X1 U1606 ( .A(n4006), .B(DATAIN[7]), .S(n186), .Z(n2769) );
  MUX2_X1 U1607 ( .A(n4005), .B(DATAIN[6]), .S(n186), .Z(n2768) );
  MUX2_X1 U1608 ( .A(n4004), .B(DATAIN[5]), .S(n186), .Z(n2767) );
  MUX2_X1 U1609 ( .A(n4003), .B(DATAIN[4]), .S(n186), .Z(n2766) );
  MUX2_X1 U1610 ( .A(n4002), .B(DATAIN[3]), .S(n186), .Z(n2765) );
  MUX2_X1 U1611 ( .A(n4001), .B(DATAIN[2]), .S(n186), .Z(n2764) );
  MUX2_X1 U1612 ( .A(n4000), .B(DATAIN[1]), .S(n186), .Z(n2763) );
  MUX2_X1 U1613 ( .A(n3999), .B(DATAIN[0]), .S(n186), .Z(n2762) );
  AND2_X1 U1614 ( .A1(n1184), .A2(n763), .ZN(n1185) );
  NOR3_X1 U1615 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n1186), .ZN(n763) );
  MUX2_X1 U1616 ( .A(n1187), .B(DATAIN[31]), .S(n191), .Z(n2761) );
  MUX2_X1 U1617 ( .A(n1189), .B(DATAIN[30]), .S(n191), .Z(n2760) );
  MUX2_X1 U1618 ( .A(n1190), .B(DATAIN[29]), .S(n191), .Z(n2759) );
  MUX2_X1 U1619 ( .A(n1191), .B(DATAIN[28]), .S(n191), .Z(n2758) );
  MUX2_X1 U1620 ( .A(n1192), .B(DATAIN[27]), .S(n191), .Z(n2757) );
  MUX2_X1 U1621 ( .A(n1193), .B(DATAIN[26]), .S(n191), .Z(n2756) );
  MUX2_X1 U1622 ( .A(n1194), .B(DATAIN[25]), .S(n191), .Z(n2755) );
  MUX2_X1 U1623 ( .A(n1195), .B(DATAIN[24]), .S(n191), .Z(n2754) );
  MUX2_X1 U1624 ( .A(n1196), .B(DATAIN[23]), .S(n190), .Z(n2753) );
  MUX2_X1 U1625 ( .A(n1197), .B(DATAIN[22]), .S(n190), .Z(n2752) );
  MUX2_X1 U1626 ( .A(n1198), .B(DATAIN[21]), .S(n190), .Z(n2751) );
  MUX2_X1 U1627 ( .A(n1199), .B(DATAIN[20]), .S(n190), .Z(n2750) );
  MUX2_X1 U1628 ( .A(n1200), .B(DATAIN[19]), .S(n190), .Z(n2749) );
  MUX2_X1 U1629 ( .A(n1201), .B(DATAIN[18]), .S(n190), .Z(n2748) );
  MUX2_X1 U1630 ( .A(n1202), .B(DATAIN[17]), .S(n190), .Z(n2747) );
  MUX2_X1 U1631 ( .A(n1203), .B(DATAIN[16]), .S(n190), .Z(n2746) );
  MUX2_X1 U1632 ( .A(n1204), .B(DATAIN[15]), .S(n190), .Z(n2745) );
  MUX2_X1 U1633 ( .A(n1205), .B(DATAIN[14]), .S(n190), .Z(n2744) );
  MUX2_X1 U1634 ( .A(n1206), .B(DATAIN[13]), .S(n190), .Z(n2743) );
  MUX2_X1 U1635 ( .A(n1207), .B(DATAIN[12]), .S(n190), .Z(n2742) );
  MUX2_X1 U1636 ( .A(n1208), .B(DATAIN[11]), .S(n189), .Z(n2741) );
  MUX2_X1 U1637 ( .A(n1209), .B(DATAIN[10]), .S(n189), .Z(n2740) );
  MUX2_X1 U1638 ( .A(n1210), .B(DATAIN[9]), .S(n189), .Z(n2739) );
  MUX2_X1 U1639 ( .A(n1211), .B(DATAIN[8]), .S(n189), .Z(n2738) );
  MUX2_X1 U1640 ( .A(n1212), .B(DATAIN[7]), .S(n189), .Z(n2737) );
  MUX2_X1 U1641 ( .A(n1213), .B(DATAIN[6]), .S(n189), .Z(n2736) );
  MUX2_X1 U1642 ( .A(n1214), .B(DATAIN[5]), .S(n189), .Z(n2735) );
  MUX2_X1 U1643 ( .A(n1215), .B(DATAIN[4]), .S(n189), .Z(n2734) );
  MUX2_X1 U1644 ( .A(n1216), .B(DATAIN[3]), .S(n189), .Z(n2733) );
  MUX2_X1 U1645 ( .A(n1217), .B(DATAIN[2]), .S(n189), .Z(n2732) );
  MUX2_X1 U1646 ( .A(n1218), .B(DATAIN[1]), .S(n189), .Z(n2731) );
  MUX2_X1 U1647 ( .A(n1219), .B(DATAIN[0]), .S(n189), .Z(n2730) );
  AND2_X1 U1648 ( .A1(n1184), .A2(n766), .ZN(n1188) );
  NOR3_X1 U1649 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n1220), .ZN(n766) );
  INV_X1 U1650 ( .A(n1221), .ZN(n2729) );
  MUX2_X1 U1651 ( .A(n837), .B(n593), .S(n194), .Z(n1221) );
  INV_X1 U1652 ( .A(n1223), .ZN(n2728) );
  MUX2_X1 U1653 ( .A(n838), .B(n592), .S(n194), .Z(n1223) );
  INV_X1 U1654 ( .A(n1224), .ZN(n2727) );
  MUX2_X1 U1655 ( .A(n839), .B(n591), .S(n194), .Z(n1224) );
  INV_X1 U1656 ( .A(n1225), .ZN(n2726) );
  MUX2_X1 U1657 ( .A(n840), .B(n590), .S(n194), .Z(n1225) );
  INV_X1 U1658 ( .A(n1226), .ZN(n2725) );
  MUX2_X1 U1659 ( .A(n841), .B(n589), .S(n194), .Z(n1226) );
  INV_X1 U1660 ( .A(n1227), .ZN(n2724) );
  MUX2_X1 U1661 ( .A(n842), .B(n588), .S(n194), .Z(n1227) );
  INV_X1 U1662 ( .A(n1228), .ZN(n2723) );
  MUX2_X1 U1663 ( .A(n843), .B(n587), .S(n194), .Z(n1228) );
  INV_X1 U1664 ( .A(n1229), .ZN(n2722) );
  MUX2_X1 U1665 ( .A(n844), .B(n586), .S(n194), .Z(n1229) );
  INV_X1 U1666 ( .A(n1230), .ZN(n2721) );
  MUX2_X1 U1667 ( .A(n845), .B(n585), .S(n193), .Z(n1230) );
  INV_X1 U1668 ( .A(n1231), .ZN(n2720) );
  MUX2_X1 U1669 ( .A(n846), .B(n584), .S(n193), .Z(n1231) );
  INV_X1 U1670 ( .A(n1232), .ZN(n2719) );
  MUX2_X1 U1671 ( .A(n847), .B(n583), .S(n193), .Z(n1232) );
  INV_X1 U1672 ( .A(n1233), .ZN(n2718) );
  MUX2_X1 U1673 ( .A(n848), .B(n582), .S(n193), .Z(n1233) );
  INV_X1 U1674 ( .A(n1234), .ZN(n2717) );
  MUX2_X1 U1675 ( .A(n849), .B(n581), .S(n193), .Z(n1234) );
  INV_X1 U1676 ( .A(n1235), .ZN(n2716) );
  MUX2_X1 U1677 ( .A(n850), .B(n580), .S(n193), .Z(n1235) );
  INV_X1 U1678 ( .A(n1236), .ZN(n2715) );
  MUX2_X1 U1679 ( .A(n851), .B(n579), .S(n193), .Z(n1236) );
  INV_X1 U1680 ( .A(n1237), .ZN(n2714) );
  MUX2_X1 U1681 ( .A(n852), .B(n578), .S(n193), .Z(n1237) );
  INV_X1 U1682 ( .A(n1238), .ZN(n2713) );
  MUX2_X1 U1683 ( .A(n853), .B(n577), .S(n193), .Z(n1238) );
  INV_X1 U1684 ( .A(n1239), .ZN(n2712) );
  MUX2_X1 U1685 ( .A(n854), .B(n576), .S(n193), .Z(n1239) );
  INV_X1 U1686 ( .A(n1240), .ZN(n2711) );
  MUX2_X1 U1687 ( .A(n855), .B(n575), .S(n193), .Z(n1240) );
  INV_X1 U1688 ( .A(n1241), .ZN(n2710) );
  MUX2_X1 U1689 ( .A(n856), .B(n574), .S(n193), .Z(n1241) );
  INV_X1 U1690 ( .A(n1242), .ZN(n2709) );
  MUX2_X1 U1691 ( .A(n857), .B(n573), .S(n192), .Z(n1242) );
  INV_X1 U1692 ( .A(n1243), .ZN(n2708) );
  MUX2_X1 U1693 ( .A(n858), .B(n572), .S(n192), .Z(n1243) );
  INV_X1 U1694 ( .A(n1244), .ZN(n2707) );
  MUX2_X1 U1695 ( .A(n859), .B(n571), .S(n192), .Z(n1244) );
  INV_X1 U1696 ( .A(n1245), .ZN(n2706) );
  MUX2_X1 U1697 ( .A(n860), .B(n570), .S(n192), .Z(n1245) );
  INV_X1 U1698 ( .A(n1246), .ZN(n2705) );
  MUX2_X1 U1699 ( .A(n861), .B(n569), .S(n192), .Z(n1246) );
  INV_X1 U1700 ( .A(n1247), .ZN(n2704) );
  MUX2_X1 U1701 ( .A(n862), .B(n568), .S(n192), .Z(n1247) );
  INV_X1 U1702 ( .A(n1248), .ZN(n2703) );
  MUX2_X1 U1703 ( .A(n863), .B(n567), .S(n192), .Z(n1248) );
  INV_X1 U1704 ( .A(n1249), .ZN(n2702) );
  MUX2_X1 U1705 ( .A(n864), .B(n566), .S(n192), .Z(n1249) );
  INV_X1 U1706 ( .A(n1250), .ZN(n2701) );
  MUX2_X1 U1707 ( .A(n865), .B(n565), .S(n192), .Z(n1250) );
  INV_X1 U1708 ( .A(n1251), .ZN(n2700) );
  MUX2_X1 U1709 ( .A(n866), .B(n564), .S(n192), .Z(n1251) );
  INV_X1 U1710 ( .A(n1252), .ZN(n2699) );
  MUX2_X1 U1711 ( .A(n867), .B(n563), .S(n192), .Z(n1252) );
  INV_X1 U1712 ( .A(n1253), .ZN(n2698) );
  MUX2_X1 U1713 ( .A(n868), .B(n562), .S(n192), .Z(n1253) );
  AND2_X1 U1714 ( .A1(n1184), .A2(n768), .ZN(n1222) );
  NOR3_X1 U1715 ( .A1(n1186), .A2(ADD_WR[2]), .A3(n1220), .ZN(n768) );
  MUX2_X1 U1716 ( .A(n3998), .B(DATAIN[31]), .S(n197), .Z(n2697) );
  MUX2_X1 U1717 ( .A(n3997), .B(DATAIN[30]), .S(n197), .Z(n2696) );
  MUX2_X1 U1718 ( .A(n3996), .B(DATAIN[29]), .S(n197), .Z(n2695) );
  MUX2_X1 U1719 ( .A(n3995), .B(DATAIN[28]), .S(n197), .Z(n2694) );
  MUX2_X1 U1720 ( .A(n3994), .B(DATAIN[27]), .S(n197), .Z(n2693) );
  MUX2_X1 U1721 ( .A(n3993), .B(DATAIN[26]), .S(n197), .Z(n2692) );
  MUX2_X1 U1722 ( .A(n3992), .B(DATAIN[25]), .S(n197), .Z(n2691) );
  MUX2_X1 U1723 ( .A(n3991), .B(DATAIN[24]), .S(n197), .Z(n2690) );
  MUX2_X1 U1724 ( .A(n3990), .B(DATAIN[23]), .S(n196), .Z(n2689) );
  MUX2_X1 U1725 ( .A(n3989), .B(DATAIN[22]), .S(n196), .Z(n2688) );
  MUX2_X1 U1726 ( .A(n3988), .B(DATAIN[21]), .S(n196), .Z(n2687) );
  MUX2_X1 U1727 ( .A(n3987), .B(DATAIN[20]), .S(n196), .Z(n2686) );
  MUX2_X1 U1728 ( .A(n3986), .B(DATAIN[19]), .S(n196), .Z(n2685) );
  MUX2_X1 U1729 ( .A(n3985), .B(DATAIN[18]), .S(n196), .Z(n2684) );
  MUX2_X1 U1730 ( .A(n3984), .B(DATAIN[17]), .S(n196), .Z(n2683) );
  MUX2_X1 U1731 ( .A(n3983), .B(DATAIN[16]), .S(n196), .Z(n2682) );
  MUX2_X1 U1732 ( .A(n3982), .B(DATAIN[15]), .S(n196), .Z(n2681) );
  MUX2_X1 U1733 ( .A(n3981), .B(DATAIN[14]), .S(n196), .Z(n2680) );
  MUX2_X1 U1734 ( .A(n3980), .B(DATAIN[13]), .S(n196), .Z(n2679) );
  MUX2_X1 U1735 ( .A(n3979), .B(DATAIN[12]), .S(n196), .Z(n2678) );
  MUX2_X1 U1736 ( .A(n3978), .B(DATAIN[11]), .S(n195), .Z(n2677) );
  MUX2_X1 U1737 ( .A(n3977), .B(DATAIN[10]), .S(n195), .Z(n2676) );
  MUX2_X1 U1738 ( .A(n3976), .B(DATAIN[9]), .S(n195), .Z(n2675) );
  MUX2_X1 U1739 ( .A(n3975), .B(DATAIN[8]), .S(n195), .Z(n2674) );
  MUX2_X1 U1740 ( .A(n3974), .B(DATAIN[7]), .S(n195), .Z(n2673) );
  MUX2_X1 U1741 ( .A(n3973), .B(DATAIN[6]), .S(n195), .Z(n2672) );
  MUX2_X1 U1742 ( .A(n3972), .B(DATAIN[5]), .S(n195), .Z(n2671) );
  MUX2_X1 U1743 ( .A(n3971), .B(DATAIN[4]), .S(n195), .Z(n2670) );
  MUX2_X1 U1744 ( .A(n3970), .B(DATAIN[3]), .S(n195), .Z(n2669) );
  MUX2_X1 U1745 ( .A(n3969), .B(DATAIN[2]), .S(n195), .Z(n2668) );
  MUX2_X1 U1746 ( .A(n3968), .B(DATAIN[1]), .S(n195), .Z(n2667) );
  MUX2_X1 U1747 ( .A(n3967), .B(DATAIN[0]), .S(n195), .Z(n2666) );
  AND2_X1 U1748 ( .A1(n1184), .A2(n802), .ZN(n1254) );
  AND3_X1 U1749 ( .A1(n1186), .A2(n1220), .A3(ADD_WR[2]), .ZN(n802) );
  MUX2_X1 U1750 ( .A(n3966), .B(DATAIN[31]), .S(n200), .Z(n2665) );
  MUX2_X1 U1751 ( .A(n3965), .B(DATAIN[30]), .S(n200), .Z(n2664) );
  MUX2_X1 U1752 ( .A(n3964), .B(DATAIN[29]), .S(n200), .Z(n2663) );
  MUX2_X1 U1753 ( .A(n3963), .B(DATAIN[28]), .S(n200), .Z(n2662) );
  MUX2_X1 U1754 ( .A(n3962), .B(DATAIN[27]), .S(n200), .Z(n2661) );
  MUX2_X1 U1755 ( .A(n3961), .B(DATAIN[26]), .S(n200), .Z(n2660) );
  MUX2_X1 U1756 ( .A(n3960), .B(DATAIN[25]), .S(n200), .Z(n2659) );
  MUX2_X1 U1757 ( .A(n3959), .B(DATAIN[24]), .S(n200), .Z(n2658) );
  MUX2_X1 U1758 ( .A(n3958), .B(DATAIN[23]), .S(n199), .Z(n2657) );
  MUX2_X1 U1759 ( .A(n3957), .B(DATAIN[22]), .S(n199), .Z(n2656) );
  MUX2_X1 U1760 ( .A(n3956), .B(DATAIN[21]), .S(n199), .Z(n2655) );
  MUX2_X1 U1761 ( .A(n3955), .B(DATAIN[20]), .S(n199), .Z(n2654) );
  MUX2_X1 U1762 ( .A(n3954), .B(DATAIN[19]), .S(n199), .Z(n2653) );
  MUX2_X1 U1763 ( .A(n3953), .B(DATAIN[18]), .S(n199), .Z(n2652) );
  MUX2_X1 U1764 ( .A(n3952), .B(DATAIN[17]), .S(n199), .Z(n2651) );
  MUX2_X1 U1765 ( .A(n3951), .B(DATAIN[16]), .S(n199), .Z(n2650) );
  MUX2_X1 U1766 ( .A(n3950), .B(DATAIN[15]), .S(n199), .Z(n2649) );
  MUX2_X1 U1767 ( .A(n3949), .B(DATAIN[14]), .S(n199), .Z(n2648) );
  MUX2_X1 U1768 ( .A(n3948), .B(DATAIN[13]), .S(n199), .Z(n2647) );
  MUX2_X1 U1769 ( .A(n3947), .B(DATAIN[12]), .S(n199), .Z(n2646) );
  MUX2_X1 U1770 ( .A(n3946), .B(DATAIN[11]), .S(n198), .Z(n2645) );
  MUX2_X1 U1771 ( .A(n3945), .B(DATAIN[10]), .S(n198), .Z(n2644) );
  MUX2_X1 U1772 ( .A(n3944), .B(DATAIN[9]), .S(n198), .Z(n2643) );
  MUX2_X1 U1773 ( .A(n3943), .B(DATAIN[8]), .S(n198), .Z(n2642) );
  MUX2_X1 U1774 ( .A(n3942), .B(DATAIN[7]), .S(n198), .Z(n2641) );
  MUX2_X1 U1775 ( .A(n3941), .B(DATAIN[6]), .S(n198), .Z(n2640) );
  MUX2_X1 U1776 ( .A(n3940), .B(DATAIN[5]), .S(n198), .Z(n2639) );
  MUX2_X1 U1777 ( .A(n3939), .B(DATAIN[4]), .S(n198), .Z(n2638) );
  MUX2_X1 U1778 ( .A(n3938), .B(DATAIN[3]), .S(n198), .Z(n2637) );
  MUX2_X1 U1779 ( .A(n3937), .B(DATAIN[2]), .S(n198), .Z(n2636) );
  MUX2_X1 U1780 ( .A(n3936), .B(DATAIN[1]), .S(n198), .Z(n2635) );
  MUX2_X1 U1781 ( .A(n3935), .B(DATAIN[0]), .S(n198), .Z(n2634) );
  AND2_X1 U1782 ( .A1(n1184), .A2(n836), .ZN(n1255) );
  AND3_X1 U1783 ( .A1(ADD_WR[0]), .A2(n1220), .A3(ADD_WR[2]), .ZN(n836) );
  INV_X1 U1784 ( .A(n1256), .ZN(n2633) );
  MUX2_X1 U1785 ( .A(n933), .B(n593), .S(n203), .Z(n1256) );
  INV_X1 U1786 ( .A(n1258), .ZN(n2632) );
  MUX2_X1 U1787 ( .A(n934), .B(n592), .S(n203), .Z(n1258) );
  INV_X1 U1788 ( .A(n1259), .ZN(n2631) );
  MUX2_X1 U1789 ( .A(n935), .B(n591), .S(n203), .Z(n1259) );
  INV_X1 U1790 ( .A(n1260), .ZN(n2630) );
  MUX2_X1 U1791 ( .A(n936), .B(n590), .S(n203), .Z(n1260) );
  INV_X1 U1792 ( .A(n1261), .ZN(n2629) );
  MUX2_X1 U1793 ( .A(n937), .B(n589), .S(n203), .Z(n1261) );
  INV_X1 U1794 ( .A(n1262), .ZN(n2628) );
  MUX2_X1 U1795 ( .A(n938), .B(n588), .S(n203), .Z(n1262) );
  INV_X1 U1796 ( .A(n1263), .ZN(n2627) );
  MUX2_X1 U1797 ( .A(n939), .B(n587), .S(n203), .Z(n1263) );
  INV_X1 U1798 ( .A(n1264), .ZN(n2626) );
  MUX2_X1 U1799 ( .A(n940), .B(n586), .S(n203), .Z(n1264) );
  INV_X1 U1800 ( .A(n1265), .ZN(n2625) );
  MUX2_X1 U1801 ( .A(n941), .B(n585), .S(n202), .Z(n1265) );
  INV_X1 U1802 ( .A(n1266), .ZN(n2624) );
  MUX2_X1 U1803 ( .A(n942), .B(n584), .S(n202), .Z(n1266) );
  INV_X1 U1804 ( .A(n1267), .ZN(n2623) );
  MUX2_X1 U1805 ( .A(n943), .B(n583), .S(n202), .Z(n1267) );
  INV_X1 U1806 ( .A(n1268), .ZN(n2622) );
  MUX2_X1 U1807 ( .A(n944), .B(n582), .S(n202), .Z(n1268) );
  INV_X1 U1808 ( .A(n1269), .ZN(n2621) );
  MUX2_X1 U1809 ( .A(n945), .B(n581), .S(n202), .Z(n1269) );
  INV_X1 U1810 ( .A(n1270), .ZN(n2620) );
  MUX2_X1 U1811 ( .A(n946), .B(n580), .S(n202), .Z(n1270) );
  INV_X1 U1812 ( .A(n1271), .ZN(n2619) );
  MUX2_X1 U1813 ( .A(n947), .B(n579), .S(n202), .Z(n1271) );
  INV_X1 U1814 ( .A(n1272), .ZN(n2618) );
  MUX2_X1 U1815 ( .A(n948), .B(n578), .S(n202), .Z(n1272) );
  INV_X1 U1816 ( .A(n1273), .ZN(n2617) );
  MUX2_X1 U1817 ( .A(n949), .B(n577), .S(n202), .Z(n1273) );
  INV_X1 U1818 ( .A(n1274), .ZN(n2616) );
  MUX2_X1 U1819 ( .A(n950), .B(n576), .S(n202), .Z(n1274) );
  INV_X1 U1820 ( .A(n1275), .ZN(n2615) );
  MUX2_X1 U1821 ( .A(n951), .B(n575), .S(n202), .Z(n1275) );
  INV_X1 U1822 ( .A(n1276), .ZN(n2614) );
  MUX2_X1 U1823 ( .A(n952), .B(n574), .S(n202), .Z(n1276) );
  INV_X1 U1824 ( .A(n1277), .ZN(n2613) );
  MUX2_X1 U1825 ( .A(n953), .B(n573), .S(n201), .Z(n1277) );
  INV_X1 U1826 ( .A(n1278), .ZN(n2612) );
  MUX2_X1 U1827 ( .A(n954), .B(n572), .S(n201), .Z(n1278) );
  INV_X1 U1828 ( .A(n1279), .ZN(n2611) );
  MUX2_X1 U1829 ( .A(n955), .B(n571), .S(n201), .Z(n1279) );
  INV_X1 U1830 ( .A(n1280), .ZN(n2610) );
  MUX2_X1 U1831 ( .A(n956), .B(n570), .S(n201), .Z(n1280) );
  INV_X1 U1832 ( .A(n1281), .ZN(n2609) );
  MUX2_X1 U1833 ( .A(n957), .B(n569), .S(n201), .Z(n1281) );
  INV_X1 U1834 ( .A(n1282), .ZN(n2608) );
  MUX2_X1 U1835 ( .A(n958), .B(n568), .S(n201), .Z(n1282) );
  INV_X1 U1836 ( .A(n1283), .ZN(n2607) );
  MUX2_X1 U1837 ( .A(n959), .B(n567), .S(n201), .Z(n1283) );
  INV_X1 U1838 ( .A(n1284), .ZN(n2606) );
  MUX2_X1 U1839 ( .A(n960), .B(n566), .S(n201), .Z(n1284) );
  INV_X1 U1840 ( .A(n1285), .ZN(n2605) );
  MUX2_X1 U1841 ( .A(n961), .B(n565), .S(n201), .Z(n1285) );
  INV_X1 U1842 ( .A(n1286), .ZN(n2604) );
  MUX2_X1 U1843 ( .A(n962), .B(n564), .S(n201), .Z(n1286) );
  INV_X1 U1844 ( .A(n1287), .ZN(n2603) );
  MUX2_X1 U1845 ( .A(n963), .B(n563), .S(n201), .Z(n1287) );
  INV_X1 U1846 ( .A(n1288), .ZN(n2602) );
  MUX2_X1 U1847 ( .A(n964), .B(n562), .S(n201), .Z(n1288) );
  AND2_X1 U1848 ( .A1(n1184), .A2(n870), .ZN(n1257) );
  AND3_X1 U1849 ( .A1(ADD_WR[1]), .A2(n1186), .A3(ADD_WR[2]), .ZN(n870) );
  MUX2_X1 U1850 ( .A(n1289), .B(DATAIN[31]), .S(n206), .Z(n2601) );
  MUX2_X1 U1851 ( .A(n1291), .B(DATAIN[30]), .S(n206), .Z(n2600) );
  MUX2_X1 U1852 ( .A(n1292), .B(DATAIN[29]), .S(n206), .Z(n2599) );
  MUX2_X1 U1853 ( .A(n1293), .B(DATAIN[28]), .S(n206), .Z(n2598) );
  MUX2_X1 U1854 ( .A(n1294), .B(DATAIN[27]), .S(n206), .Z(n2597) );
  MUX2_X1 U1855 ( .A(n1295), .B(DATAIN[26]), .S(n206), .Z(n2596) );
  MUX2_X1 U1856 ( .A(n1296), .B(DATAIN[25]), .S(n206), .Z(n2595) );
  MUX2_X1 U1857 ( .A(n1297), .B(DATAIN[24]), .S(n206), .Z(n2594) );
  MUX2_X1 U1858 ( .A(n1298), .B(DATAIN[23]), .S(n205), .Z(n2593) );
  MUX2_X1 U1859 ( .A(n1299), .B(DATAIN[22]), .S(n205), .Z(n2592) );
  MUX2_X1 U1860 ( .A(n1300), .B(DATAIN[21]), .S(n205), .Z(n2591) );
  MUX2_X1 U1861 ( .A(n1301), .B(DATAIN[20]), .S(n205), .Z(n2590) );
  MUX2_X1 U1862 ( .A(n1302), .B(DATAIN[19]), .S(n205), .Z(n2589) );
  MUX2_X1 U1863 ( .A(n1303), .B(DATAIN[18]), .S(n205), .Z(n2588) );
  MUX2_X1 U1864 ( .A(n1304), .B(DATAIN[17]), .S(n205), .Z(n2587) );
  MUX2_X1 U1865 ( .A(n1305), .B(DATAIN[16]), .S(n205), .Z(n2586) );
  MUX2_X1 U1866 ( .A(n1306), .B(DATAIN[15]), .S(n205), .Z(n2585) );
  MUX2_X1 U1867 ( .A(n1307), .B(DATAIN[14]), .S(n205), .Z(n2584) );
  MUX2_X1 U1868 ( .A(n1308), .B(DATAIN[13]), .S(n205), .Z(n2583) );
  MUX2_X1 U1869 ( .A(n1309), .B(DATAIN[12]), .S(n205), .Z(n2582) );
  MUX2_X1 U1870 ( .A(n1310), .B(DATAIN[11]), .S(n204), .Z(n2581) );
  MUX2_X1 U1871 ( .A(n1311), .B(DATAIN[10]), .S(n204), .Z(n2580) );
  MUX2_X1 U1872 ( .A(n1312), .B(DATAIN[9]), .S(n204), .Z(n2579) );
  MUX2_X1 U1873 ( .A(n1313), .B(DATAIN[8]), .S(n204), .Z(n2578) );
  MUX2_X1 U1874 ( .A(n1314), .B(DATAIN[7]), .S(n204), .Z(n2577) );
  MUX2_X1 U1875 ( .A(n1315), .B(DATAIN[6]), .S(n204), .Z(n2576) );
  MUX2_X1 U1876 ( .A(n1316), .B(DATAIN[5]), .S(n204), .Z(n2575) );
  MUX2_X1 U1877 ( .A(n1317), .B(DATAIN[4]), .S(n204), .Z(n2574) );
  MUX2_X1 U1878 ( .A(n1318), .B(DATAIN[3]), .S(n204), .Z(n2573) );
  MUX2_X1 U1879 ( .A(n1319), .B(DATAIN[2]), .S(n204), .Z(n2572) );
  MUX2_X1 U1880 ( .A(n1320), .B(DATAIN[1]), .S(n204), .Z(n2571) );
  MUX2_X1 U1881 ( .A(n1321), .B(DATAIN[0]), .S(n204), .Z(n2570) );
  AND2_X1 U1882 ( .A1(n1184), .A2(n872), .ZN(n1290) );
  AND3_X1 U1883 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n872) );
  AND3_X1 U1884 ( .A1(ADD_WR[3]), .A2(n875), .A3(ADD_WR[4]), .ZN(n1184) );
  NOR2_X1 U1885 ( .A1(n1322), .A2(n1323), .ZN(n875) );
  INV_X1 U1886 ( .A(ENABLE), .ZN(n1322) );
  OAI222_X1 U1887 ( .A1(n593), .A2(n209), .B1(n1325), .B2(n212), .C1(n3934), 
        .C2(n215), .ZN(n2569) );
  NOR4_X1 U1888 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1325)
         );
  OAI221_X1 U1889 ( .B1(n837), .B2(n218), .C1(n1333), .C2(n221), .A(n1335), 
        .ZN(n1331) );
  AOI22_X1 U1890 ( .A1(n224), .A2(n4062), .B1(n225), .B2(n1187), .ZN(n1335) );
  OAI221_X1 U1891 ( .B1(n1338), .B2(n294), .C1(n933), .C2(n297), .A(n1341), 
        .ZN(n1330) );
  AOI22_X1 U1892 ( .A1(n300), .A2(n1289), .B1(n303), .B2(n4030), .ZN(n1341) );
  OAI211_X1 U1893 ( .C1(n517), .C2(n306), .A(n1345), .B(n1346), .ZN(n1329) );
  AOI221_X1 U1894 ( .B1(n307), .B2(n1148), .C1(n312), .C2(n4158), .A(n1349), 
        .ZN(n1346) );
  OAI22_X1 U1895 ( .A1(n613), .A2(n315), .B1(n1351), .B2(n318), .ZN(n1349) );
  AOI22_X1 U1896 ( .A1(n321), .A2(n4190), .B1(n324), .B2(n1046), .ZN(n1345) );
  NAND4_X1 U1897 ( .A1(n1358), .A2(n1356), .A3(n1357), .A4(n1355), .ZN(n1328)
         );
  AOI221_X1 U1898 ( .B1(n327), .B2(n4222), .C1(n330), .C2(n4254), .A(n1361), 
        .ZN(n1358) );
  OAI22_X1 U1899 ( .A1(n389), .A2(n333), .B1(n357), .B2(n20), .ZN(n1361) );
  AOI221_X1 U1900 ( .B1(n336), .B2(n4286), .C1(n339), .C2(n4318), .A(n1366), 
        .ZN(n1357) );
  OAI22_X1 U1901 ( .A1(n261), .A2(n342), .B1(n229), .B2(n343), .ZN(n1366) );
  AOI221_X1 U1902 ( .B1(n348), .B2(n769), .C1(n351), .C2(n803), .A(n1371), 
        .ZN(n1356) );
  OAI22_X1 U1903 ( .A1(n1372), .A2(n354), .B1(n1374), .B2(n421), .ZN(n1371) );
  AOI221_X1 U1904 ( .B1(n423), .B2(n730), .C1(n427), .C2(n3966), .A(n1378), 
        .ZN(n1355) );
  OAI22_X1 U1905 ( .A1(n1379), .A2(n430), .B1(n1381), .B2(n22), .ZN(n1378) );
  OAI222_X1 U1906 ( .A1(n592), .A2(n209), .B1(n1383), .B2(n212), .C1(n3933), 
        .C2(n215), .ZN(n2568) );
  NOR4_X1 U1907 ( .A1(n1384), .A2(n1385), .A3(n1386), .A4(n1387), .ZN(n1383)
         );
  OAI221_X1 U1908 ( .B1(n838), .B2(n218), .C1(n1388), .C2(n221), .A(n1389), 
        .ZN(n1387) );
  AOI22_X1 U1909 ( .A1(n224), .A2(n4061), .B1(n30), .B2(n1189), .ZN(n1389) );
  OAI221_X1 U1910 ( .B1(n1390), .B2(n294), .C1(n934), .C2(n297), .A(n1391), 
        .ZN(n1386) );
  AOI22_X1 U1911 ( .A1(n300), .A2(n1291), .B1(n303), .B2(n4029), .ZN(n1391) );
  OAI211_X1 U1912 ( .C1(n518), .C2(n306), .A(n1392), .B(n1393), .ZN(n1385) );
  AOI221_X1 U1913 ( .B1(n307), .B2(n1150), .C1(n312), .C2(n4157), .A(n1394), 
        .ZN(n1393) );
  OAI22_X1 U1914 ( .A1(n614), .A2(n315), .B1(n1395), .B2(n318), .ZN(n1394) );
  AOI22_X1 U1915 ( .A1(n321), .A2(n4189), .B1(n324), .B2(n1048), .ZN(n1392) );
  NAND4_X1 U1916 ( .A1(n1396), .A2(n1397), .A3(n1398), .A4(n1399), .ZN(n1384)
         );
  AOI221_X1 U1917 ( .B1(n327), .B2(n4221), .C1(n330), .C2(n4253), .A(n1400), 
        .ZN(n1399) );
  OAI22_X1 U1918 ( .A1(n390), .A2(n32), .B1(n358), .B2(n21), .ZN(n1400) );
  AOI221_X1 U1919 ( .B1(n336), .B2(n4285), .C1(n339), .C2(n4317), .A(n1401), 
        .ZN(n1398) );
  OAI22_X1 U1920 ( .A1(n262), .A2(n33), .B1(n230), .B2(n345), .ZN(n1401) );
  AOI221_X1 U1921 ( .B1(n348), .B2(n771), .C1(n351), .C2(n805), .A(n1402), 
        .ZN(n1397) );
  OAI22_X1 U1922 ( .A1(n1403), .A2(n354), .B1(n1404), .B2(n421), .ZN(n1402) );
  AOI221_X1 U1923 ( .B1(n423), .B2(n732), .C1(n427), .C2(n3965), .A(n1405), 
        .ZN(n1396) );
  OAI22_X1 U1924 ( .A1(n1406), .A2(n430), .B1(n1407), .B2(n5), .ZN(n1405) );
  OAI222_X1 U1925 ( .A1(n591), .A2(n209), .B1(n1408), .B2(n212), .C1(n3932), 
        .C2(n215), .ZN(n2567) );
  NOR4_X1 U1926 ( .A1(n1409), .A2(n1410), .A3(n1411), .A4(n1412), .ZN(n1408)
         );
  OAI221_X1 U1927 ( .B1(n839), .B2(n218), .C1(n1413), .C2(n221), .A(n1414), 
        .ZN(n1412) );
  AOI22_X1 U1928 ( .A1(n224), .A2(n4060), .B1(n29), .B2(n1190), .ZN(n1414) );
  OAI221_X1 U1929 ( .B1(n1415), .B2(n294), .C1(n935), .C2(n297), .A(n1416), 
        .ZN(n1411) );
  AOI22_X1 U1930 ( .A1(n300), .A2(n1292), .B1(n303), .B2(n4028), .ZN(n1416) );
  OAI211_X1 U1931 ( .C1(n519), .C2(n306), .A(n1417), .B(n1418), .ZN(n1410) );
  AOI221_X1 U1932 ( .B1(n309), .B2(n1151), .C1(n312), .C2(n4156), .A(n1419), 
        .ZN(n1418) );
  OAI22_X1 U1933 ( .A1(n615), .A2(n315), .B1(n1420), .B2(n318), .ZN(n1419) );
  AOI22_X1 U1934 ( .A1(n321), .A2(n4188), .B1(n324), .B2(n1049), .ZN(n1417) );
  NAND4_X1 U1935 ( .A1(n1424), .A2(n1422), .A3(n1423), .A4(n1421), .ZN(n1409)
         );
  AOI221_X1 U1936 ( .B1(n327), .B2(n4220), .C1(n330), .C2(n4252), .A(n1425), 
        .ZN(n1424) );
  OAI22_X1 U1937 ( .A1(n391), .A2(n332), .B1(n359), .B2(n21), .ZN(n1425) );
  AOI221_X1 U1938 ( .B1(n336), .B2(n4284), .C1(n339), .C2(n4316), .A(n1426), 
        .ZN(n1423) );
  OAI22_X1 U1939 ( .A1(n263), .A2(n34), .B1(n231), .B2(n343), .ZN(n1426) );
  AOI221_X1 U1940 ( .B1(n348), .B2(n772), .C1(n351), .C2(n806), .A(n1427), 
        .ZN(n1422) );
  OAI22_X1 U1941 ( .A1(n1428), .A2(n354), .B1(n1429), .B2(n421), .ZN(n1427) );
  AOI221_X1 U1942 ( .B1(n423), .B2(n733), .C1(n427), .C2(n3964), .A(n1430), 
        .ZN(n1421) );
  OAI22_X1 U1943 ( .A1(n1431), .A2(n430), .B1(n1432), .B2(n5), .ZN(n1430) );
  OAI222_X1 U1944 ( .A1(n590), .A2(n209), .B1(n1433), .B2(n212), .C1(n3931), 
        .C2(n215), .ZN(n2566) );
  NOR4_X1 U1945 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1433)
         );
  OAI221_X1 U1946 ( .B1(n840), .B2(n218), .C1(n1438), .C2(n221), .A(n1439), 
        .ZN(n1437) );
  AOI22_X1 U1947 ( .A1(n224), .A2(n4059), .B1(n227), .B2(n1191), .ZN(n1439) );
  OAI221_X1 U1948 ( .B1(n1440), .B2(n294), .C1(n936), .C2(n297), .A(n1441), 
        .ZN(n1436) );
  AOI22_X1 U1949 ( .A1(n300), .A2(n1293), .B1(n303), .B2(n4027), .ZN(n1441) );
  OAI211_X1 U1950 ( .C1(n520), .C2(n306), .A(n1442), .B(n1443), .ZN(n1435) );
  AOI221_X1 U1951 ( .B1(n308), .B2(n1152), .C1(n312), .C2(n4155), .A(n1444), 
        .ZN(n1443) );
  OAI22_X1 U1952 ( .A1(n616), .A2(n315), .B1(n1445), .B2(n318), .ZN(n1444) );
  AOI22_X1 U1953 ( .A1(n321), .A2(n4187), .B1(n324), .B2(n1050), .ZN(n1442) );
  NAND4_X1 U1954 ( .A1(n1449), .A2(n1447), .A3(n1448), .A4(n1446), .ZN(n1434)
         );
  AOI221_X1 U1955 ( .B1(n327), .B2(n4219), .C1(n330), .C2(n4251), .A(n1450), 
        .ZN(n1449) );
  OAI22_X1 U1956 ( .A1(n392), .A2(n31), .B1(n360), .B2(n20), .ZN(n1450) );
  AOI221_X1 U1957 ( .B1(n336), .B2(n4283), .C1(n339), .C2(n4315), .A(n1451), 
        .ZN(n1448) );
  OAI22_X1 U1958 ( .A1(n264), .A2(n341), .B1(n232), .B2(n343), .ZN(n1451) );
  AOI221_X1 U1959 ( .B1(n348), .B2(n773), .C1(n351), .C2(n807), .A(n1452), 
        .ZN(n1447) );
  OAI22_X1 U1960 ( .A1(n1453), .A2(n354), .B1(n1454), .B2(n421), .ZN(n1452) );
  AOI221_X1 U1961 ( .B1(n422), .B2(n734), .C1(n427), .C2(n3963), .A(n1455), 
        .ZN(n1446) );
  OAI22_X1 U1962 ( .A1(n1456), .A2(n430), .B1(n1457), .B2(n23), .ZN(n1455) );
  OAI222_X1 U1963 ( .A1(n589), .A2(n209), .B1(n1458), .B2(n212), .C1(n3930), 
        .C2(n215), .ZN(n2565) );
  NOR4_X1 U1964 ( .A1(n1459), .A2(n1460), .A3(n1461), .A4(n1462), .ZN(n1458)
         );
  OAI221_X1 U1965 ( .B1(n841), .B2(n218), .C1(n1463), .C2(n221), .A(n1464), 
        .ZN(n1462) );
  AOI22_X1 U1966 ( .A1(n224), .A2(n4058), .B1(n225), .B2(n1192), .ZN(n1464) );
  OAI221_X1 U1967 ( .B1(n1465), .B2(n294), .C1(n937), .C2(n297), .A(n1466), 
        .ZN(n1461) );
  AOI22_X1 U1968 ( .A1(n300), .A2(n1294), .B1(n303), .B2(n4026), .ZN(n1466) );
  OAI211_X1 U1969 ( .C1(n521), .C2(n306), .A(n1467), .B(n1468), .ZN(n1460) );
  AOI221_X1 U1970 ( .B1(n309), .B2(n1153), .C1(n312), .C2(n4154), .A(n1469), 
        .ZN(n1468) );
  OAI22_X1 U1971 ( .A1(n617), .A2(n315), .B1(n1470), .B2(n318), .ZN(n1469) );
  AOI22_X1 U1972 ( .A1(n321), .A2(n4186), .B1(n324), .B2(n1051), .ZN(n1467) );
  NAND4_X1 U1973 ( .A1(n1474), .A2(n1472), .A3(n1473), .A4(n1471), .ZN(n1459)
         );
  AOI221_X1 U1974 ( .B1(n327), .B2(n4218), .C1(n330), .C2(n4250), .A(n1475), 
        .ZN(n1474) );
  OAI22_X1 U1975 ( .A1(n393), .A2(n331), .B1(n361), .B2(n20), .ZN(n1475) );
  AOI221_X1 U1976 ( .B1(n336), .B2(n4282), .C1(n339), .C2(n4314), .A(n1476), 
        .ZN(n1473) );
  OAI22_X1 U1977 ( .A1(n265), .A2(n340), .B1(n233), .B2(n345), .ZN(n1476) );
  AOI221_X1 U1978 ( .B1(n348), .B2(n774), .C1(n351), .C2(n808), .A(n1477), 
        .ZN(n1472) );
  OAI22_X1 U1979 ( .A1(n1478), .A2(n354), .B1(n1479), .B2(n421), .ZN(n1477) );
  AOI221_X1 U1980 ( .B1(n423), .B2(n735), .C1(n427), .C2(n3962), .A(n1480), 
        .ZN(n1471) );
  OAI22_X1 U1981 ( .A1(n1481), .A2(n430), .B1(n1482), .B2(n23), .ZN(n1480) );
  OAI222_X1 U1982 ( .A1(n588), .A2(n209), .B1(n1483), .B2(n212), .C1(n3929), 
        .C2(n215), .ZN(n2564) );
  NOR4_X1 U1983 ( .A1(n1484), .A2(n1485), .A3(n1486), .A4(n1487), .ZN(n1483)
         );
  OAI221_X1 U1984 ( .B1(n842), .B2(n218), .C1(n1488), .C2(n221), .A(n1489), 
        .ZN(n1487) );
  AOI22_X1 U1985 ( .A1(n224), .A2(n4057), .B1(n30), .B2(n1193), .ZN(n1489) );
  OAI221_X1 U1986 ( .B1(n1490), .B2(n294), .C1(n938), .C2(n297), .A(n1491), 
        .ZN(n1486) );
  AOI22_X1 U1987 ( .A1(n300), .A2(n1295), .B1(n303), .B2(n4025), .ZN(n1491) );
  OAI211_X1 U1988 ( .C1(n522), .C2(n306), .A(n1492), .B(n1493), .ZN(n1485) );
  AOI221_X1 U1989 ( .B1(n308), .B2(n1154), .C1(n312), .C2(n4153), .A(n1494), 
        .ZN(n1493) );
  OAI22_X1 U1990 ( .A1(n618), .A2(n315), .B1(n1495), .B2(n318), .ZN(n1494) );
  AOI22_X1 U1991 ( .A1(n321), .A2(n4185), .B1(n324), .B2(n1052), .ZN(n1492) );
  NAND4_X1 U1992 ( .A1(n1499), .A2(n1497), .A3(n1498), .A4(n1496), .ZN(n1484)
         );
  AOI221_X1 U1993 ( .B1(n327), .B2(n4217), .C1(n330), .C2(n4249), .A(n1500), 
        .ZN(n1499) );
  OAI22_X1 U1994 ( .A1(n394), .A2(n333), .B1(n362), .B2(n20), .ZN(n1500) );
  AOI221_X1 U1995 ( .B1(n336), .B2(n4281), .C1(n339), .C2(n4313), .A(n1501), 
        .ZN(n1498) );
  OAI22_X1 U1996 ( .A1(n266), .A2(n342), .B1(n234), .B2(n345), .ZN(n1501) );
  AOI221_X1 U1997 ( .B1(n348), .B2(n775), .C1(n351), .C2(n809), .A(n1502), 
        .ZN(n1497) );
  OAI22_X1 U1998 ( .A1(n1503), .A2(n354), .B1(n1504), .B2(n421), .ZN(n1502) );
  AOI221_X1 U1999 ( .B1(n422), .B2(n736), .C1(n427), .C2(n3961), .A(n1505), 
        .ZN(n1496) );
  OAI22_X1 U2000 ( .A1(n1506), .A2(n430), .B1(n1507), .B2(n22), .ZN(n1505) );
  OAI222_X1 U2001 ( .A1(n587), .A2(n209), .B1(n1508), .B2(n212), .C1(n3928), 
        .C2(n215), .ZN(n2563) );
  NOR4_X1 U2002 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .ZN(n1508)
         );
  OAI221_X1 U2003 ( .B1(n843), .B2(n218), .C1(n1513), .C2(n221), .A(n1514), 
        .ZN(n1512) );
  AOI22_X1 U2004 ( .A1(n224), .A2(n4056), .B1(n29), .B2(n1194), .ZN(n1514) );
  OAI221_X1 U2005 ( .B1(n1515), .B2(n294), .C1(n939), .C2(n297), .A(n1516), 
        .ZN(n1511) );
  AOI22_X1 U2006 ( .A1(n300), .A2(n1296), .B1(n303), .B2(n4024), .ZN(n1516) );
  OAI211_X1 U2007 ( .C1(n523), .C2(n306), .A(n1517), .B(n1518), .ZN(n1510) );
  AOI221_X1 U2008 ( .B1(n309), .B2(n1155), .C1(n312), .C2(n4152), .A(n1519), 
        .ZN(n1518) );
  OAI22_X1 U2009 ( .A1(n619), .A2(n315), .B1(n1520), .B2(n318), .ZN(n1519) );
  AOI22_X1 U2010 ( .A1(n321), .A2(n4184), .B1(n324), .B2(n1053), .ZN(n1517) );
  NAND4_X1 U2011 ( .A1(n1524), .A2(n1522), .A3(n1523), .A4(n1521), .ZN(n1509)
         );
  AOI221_X1 U2012 ( .B1(n327), .B2(n4216), .C1(n330), .C2(n4248), .A(n1525), 
        .ZN(n1524) );
  OAI22_X1 U2013 ( .A1(n395), .A2(n332), .B1(n363), .B2(n21), .ZN(n1525) );
  AOI221_X1 U2014 ( .B1(n336), .B2(n4280), .C1(n339), .C2(n4312), .A(n1526), 
        .ZN(n1523) );
  OAI22_X1 U2015 ( .A1(n267), .A2(n33), .B1(n235), .B2(n343), .ZN(n1526) );
  AOI221_X1 U2016 ( .B1(n348), .B2(n776), .C1(n351), .C2(n810), .A(n1527), 
        .ZN(n1522) );
  OAI22_X1 U2017 ( .A1(n1528), .A2(n354), .B1(n1529), .B2(n421), .ZN(n1527) );
  AOI221_X1 U2018 ( .B1(n423), .B2(n737), .C1(n427), .C2(n3960), .A(n1530), 
        .ZN(n1521) );
  OAI22_X1 U2019 ( .A1(n1531), .A2(n430), .B1(n1532), .B2(n23), .ZN(n1530) );
  OAI222_X1 U2020 ( .A1(n586), .A2(n209), .B1(n1533), .B2(n212), .C1(n3927), 
        .C2(n215), .ZN(n2562) );
  NOR4_X1 U2021 ( .A1(n1534), .A2(n1535), .A3(n1536), .A4(n1537), .ZN(n1533)
         );
  OAI221_X1 U2022 ( .B1(n844), .B2(n218), .C1(n1538), .C2(n221), .A(n1539), 
        .ZN(n1537) );
  AOI22_X1 U2023 ( .A1(n224), .A2(n4055), .B1(n227), .B2(n1195), .ZN(n1539) );
  OAI221_X1 U2024 ( .B1(n1540), .B2(n294), .C1(n940), .C2(n297), .A(n1541), 
        .ZN(n1536) );
  AOI22_X1 U2025 ( .A1(n300), .A2(n1297), .B1(n303), .B2(n4023), .ZN(n1541) );
  OAI211_X1 U2026 ( .C1(n524), .C2(n306), .A(n1542), .B(n1543), .ZN(n1535) );
  AOI221_X1 U2027 ( .B1(n309), .B2(n1156), .C1(n312), .C2(n4151), .A(n1544), 
        .ZN(n1543) );
  OAI22_X1 U2028 ( .A1(n620), .A2(n315), .B1(n1545), .B2(n318), .ZN(n1544) );
  AOI22_X1 U2029 ( .A1(n321), .A2(n4183), .B1(n324), .B2(n1054), .ZN(n1542) );
  NAND4_X1 U2030 ( .A1(n1546), .A2(n1547), .A3(n1548), .A4(n1549), .ZN(n1534)
         );
  AOI221_X1 U2031 ( .B1(n327), .B2(n4215), .C1(n330), .C2(n4247), .A(n1550), 
        .ZN(n1549) );
  OAI22_X1 U2032 ( .A1(n396), .A2(n331), .B1(n364), .B2(n21), .ZN(n1550) );
  AOI221_X1 U2033 ( .B1(n336), .B2(n4279), .C1(n339), .C2(n4311), .A(n1551), 
        .ZN(n1548) );
  OAI22_X1 U2034 ( .A1(n268), .A2(n34), .B1(n236), .B2(n345), .ZN(n1551) );
  AOI221_X1 U2035 ( .B1(n348), .B2(n777), .C1(n351), .C2(n811), .A(n1552), 
        .ZN(n1547) );
  OAI22_X1 U2036 ( .A1(n1553), .A2(n354), .B1(n1554), .B2(n421), .ZN(n1552) );
  AOI221_X1 U2037 ( .B1(n422), .B2(n738), .C1(n427), .C2(n3959), .A(n1555), 
        .ZN(n1546) );
  OAI22_X1 U2038 ( .A1(n1556), .A2(n430), .B1(n1557), .B2(n22), .ZN(n1555) );
  OAI222_X1 U2039 ( .A1(n585), .A2(n208), .B1(n1558), .B2(n211), .C1(n3926), 
        .C2(n215), .ZN(n2561) );
  NOR4_X1 U2040 ( .A1(n1559), .A2(n1560), .A3(n1561), .A4(n1562), .ZN(n1558)
         );
  OAI221_X1 U2041 ( .B1(n845), .B2(n217), .C1(n1563), .C2(n220), .A(n1564), 
        .ZN(n1562) );
  AOI22_X1 U2042 ( .A1(n223), .A2(n4054), .B1(n225), .B2(n1196), .ZN(n1564) );
  OAI221_X1 U2043 ( .B1(n1565), .B2(n293), .C1(n941), .C2(n296), .A(n1566), 
        .ZN(n1561) );
  AOI22_X1 U2044 ( .A1(n299), .A2(n1298), .B1(n302), .B2(n4022), .ZN(n1566) );
  OAI211_X1 U2045 ( .C1(n525), .C2(n305), .A(n1567), .B(n1568), .ZN(n1560) );
  AOI221_X1 U2046 ( .B1(n307), .B2(n1157), .C1(n311), .C2(n4150), .A(n1569), 
        .ZN(n1568) );
  OAI22_X1 U2047 ( .A1(n621), .A2(n314), .B1(n1570), .B2(n317), .ZN(n1569) );
  AOI22_X1 U2048 ( .A1(n320), .A2(n4182), .B1(n323), .B2(n1055), .ZN(n1567) );
  NAND4_X1 U2049 ( .A1(n1574), .A2(n1571), .A3(n1572), .A4(n1573), .ZN(n1559)
         );
  AOI221_X1 U2050 ( .B1(n326), .B2(n4214), .C1(n329), .C2(n4246), .A(n1575), 
        .ZN(n1574) );
  OAI22_X1 U2051 ( .A1(n397), .A2(n31), .B1(n365), .B2(n21), .ZN(n1575) );
  AOI221_X1 U2052 ( .B1(n335), .B2(n4278), .C1(n338), .C2(n4310), .A(n1576), 
        .ZN(n1573) );
  OAI22_X1 U2053 ( .A1(n269), .A2(n341), .B1(n237), .B2(n344), .ZN(n1576) );
  AOI221_X1 U2054 ( .B1(n347), .B2(n778), .C1(n350), .C2(n812), .A(n1577), 
        .ZN(n1572) );
  OAI22_X1 U2055 ( .A1(n1578), .A2(n353), .B1(n1579), .B2(n356), .ZN(n1577) );
  OAI22_X1 U2056 ( .A1(n1581), .A2(n429), .B1(n1582), .B2(n5), .ZN(n1580) );
  OAI222_X1 U2057 ( .A1(n584), .A2(n208), .B1(n1583), .B2(n211), .C1(n3925), 
        .C2(n215), .ZN(n2560) );
  OAI221_X1 U2058 ( .B1(n846), .B2(n217), .C1(n1588), .C2(n220), .A(n1589), 
        .ZN(n1587) );
  AOI22_X1 U2059 ( .A1(n223), .A2(n4053), .B1(n29), .B2(n1197), .ZN(n1589) );
  OAI221_X1 U2060 ( .B1(n1590), .B2(n293), .C1(n942), .C2(n296), .A(n1591), 
        .ZN(n1586) );
  AOI22_X1 U2061 ( .A1(n299), .A2(n1299), .B1(n302), .B2(n4021), .ZN(n1591) );
  OAI211_X1 U2062 ( .C1(n526), .C2(n305), .A(n1592), .B(n1593), .ZN(n1585) );
  AOI221_X1 U2063 ( .B1(n308), .B2(n1158), .C1(n311), .C2(n4149), .A(n1594), 
        .ZN(n1593) );
  OAI22_X1 U2064 ( .A1(n622), .A2(n314), .B1(n1595), .B2(n317), .ZN(n1594) );
  AOI22_X1 U2065 ( .A1(n320), .A2(n4181), .B1(n323), .B2(n1056), .ZN(n1592) );
  NAND4_X1 U2066 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1584)
         );
  AOI221_X1 U2067 ( .B1(n326), .B2(n4213), .C1(n329), .C2(n4245), .A(n1600), 
        .ZN(n1599) );
  OAI22_X1 U2068 ( .A1(n398), .A2(n332), .B1(n366), .B2(n21), .ZN(n1600) );
  AOI221_X1 U2069 ( .B1(n335), .B2(n4277), .C1(n338), .C2(n4309), .A(n1601), 
        .ZN(n1598) );
  OAI22_X1 U2070 ( .A1(n270), .A2(n341), .B1(n238), .B2(n345), .ZN(n1601) );
  AOI221_X1 U2071 ( .B1(n347), .B2(n779), .C1(n350), .C2(n813), .A(n1602), 
        .ZN(n1597) );
  OAI22_X1 U2072 ( .A1(n1603), .A2(n353), .B1(n1604), .B2(n356), .ZN(n1602) );
  AOI221_X1 U2073 ( .B1(n422), .B2(n740), .C1(n426), .C2(n3957), .A(n1605), 
        .ZN(n1596) );
  OAI22_X1 U2074 ( .A1(n1606), .A2(n429), .B1(n1607), .B2(n23), .ZN(n1605) );
  OAI222_X1 U2075 ( .A1(n583), .A2(n208), .B1(n1608), .B2(n211), .C1(n3924), 
        .C2(n214), .ZN(n2559) );
  NOR4_X1 U2076 ( .A1(n1609), .A2(n1610), .A3(n1611), .A4(n1612), .ZN(n1608)
         );
  OAI221_X1 U2077 ( .B1(n847), .B2(n217), .C1(n1613), .C2(n220), .A(n1614), 
        .ZN(n1612) );
  AOI22_X1 U2078 ( .A1(n223), .A2(n4052), .B1(n30), .B2(n1198), .ZN(n1614) );
  OAI221_X1 U2079 ( .B1(n1615), .B2(n293), .C1(n943), .C2(n296), .A(n1616), 
        .ZN(n1611) );
  AOI22_X1 U2080 ( .A1(n299), .A2(n1300), .B1(n302), .B2(n4020), .ZN(n1616) );
  OAI211_X1 U2081 ( .C1(n527), .C2(n305), .A(n1617), .B(n1618), .ZN(n1610) );
  AOI221_X1 U2082 ( .B1(n307), .B2(n1159), .C1(n311), .C2(n4148), .A(n1619), 
        .ZN(n1618) );
  OAI22_X1 U2083 ( .A1(n623), .A2(n314), .B1(n1620), .B2(n317), .ZN(n1619) );
  AOI22_X1 U2084 ( .A1(n320), .A2(n4180), .B1(n323), .B2(n1057), .ZN(n1617) );
  NAND4_X1 U2085 ( .A1(n1624), .A2(n1621), .A3(n1622), .A4(n1623), .ZN(n1609)
         );
  AOI221_X1 U2086 ( .B1(n326), .B2(n4212), .C1(n329), .C2(n4244), .A(n1625), 
        .ZN(n1624) );
  OAI22_X1 U2087 ( .A1(n399), .A2(n332), .B1(n367), .B2(n20), .ZN(n1625) );
  AOI221_X1 U2088 ( .B1(n335), .B2(n4276), .C1(n338), .C2(n4308), .A(n1626), 
        .ZN(n1623) );
  OAI22_X1 U2089 ( .A1(n271), .A2(n340), .B1(n239), .B2(n344), .ZN(n1626) );
  AOI221_X1 U2090 ( .B1(n347), .B2(n780), .C1(n350), .C2(n814), .A(n1627), 
        .ZN(n1622) );
  OAI22_X1 U2091 ( .A1(n1628), .A2(n353), .B1(n1629), .B2(n356), .ZN(n1627) );
  OAI22_X1 U2092 ( .A1(n1631), .A2(n429), .B1(n1632), .B2(n23), .ZN(n1630) );
  OAI222_X1 U2093 ( .A1(n582), .A2(n208), .B1(n1633), .B2(n211), .C1(n3923), 
        .C2(n214), .ZN(n2558) );
  OAI221_X1 U2094 ( .B1(n848), .B2(n217), .C1(n1638), .C2(n220), .A(n1639), 
        .ZN(n1637) );
  AOI22_X1 U2095 ( .A1(n223), .A2(n4051), .B1(n227), .B2(n1199), .ZN(n1639) );
  OAI221_X1 U2096 ( .B1(n1640), .B2(n293), .C1(n944), .C2(n296), .A(n1641), 
        .ZN(n1636) );
  AOI22_X1 U2097 ( .A1(n299), .A2(n1301), .B1(n302), .B2(n4019), .ZN(n1641) );
  OAI211_X1 U2098 ( .C1(n528), .C2(n305), .A(n1642), .B(n1643), .ZN(n1635) );
  AOI221_X1 U2099 ( .B1(n309), .B2(n1160), .C1(n311), .C2(n4147), .A(n1644), 
        .ZN(n1643) );
  OAI22_X1 U2100 ( .A1(n624), .A2(n314), .B1(n1645), .B2(n317), .ZN(n1644) );
  AOI22_X1 U2101 ( .A1(n320), .A2(n4179), .B1(n323), .B2(n1058), .ZN(n1642) );
  NAND4_X1 U2102 ( .A1(n1646), .A2(n1647), .A3(n1648), .A4(n1649), .ZN(n1634)
         );
  AOI221_X1 U2103 ( .B1(n326), .B2(n4211), .C1(n329), .C2(n4243), .A(n1650), 
        .ZN(n1649) );
  OAI22_X1 U2104 ( .A1(n400), .A2(n333), .B1(n368), .B2(n20), .ZN(n1650) );
  AOI221_X1 U2105 ( .B1(n335), .B2(n4275), .C1(n338), .C2(n4307), .A(n1651), 
        .ZN(n1648) );
  OAI22_X1 U2106 ( .A1(n272), .A2(n340), .B1(n240), .B2(n343), .ZN(n1651) );
  AOI221_X1 U2107 ( .B1(n347), .B2(n781), .C1(n350), .C2(n815), .A(n1652), 
        .ZN(n1647) );
  OAI22_X1 U2108 ( .A1(n1653), .A2(n353), .B1(n1654), .B2(n356), .ZN(n1652) );
  AOI221_X1 U2109 ( .B1(n423), .B2(n742), .C1(n426), .C2(n3955), .A(n1655), 
        .ZN(n1646) );
  OAI22_X1 U2110 ( .A1(n1656), .A2(n429), .B1(n1657), .B2(n22), .ZN(n1655) );
  OAI222_X1 U2111 ( .A1(n581), .A2(n208), .B1(n1658), .B2(n211), .C1(n3922), 
        .C2(n214), .ZN(n2557) );
  NOR4_X1 U2112 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1658)
         );
  OAI221_X1 U2113 ( .B1(n849), .B2(n217), .C1(n1663), .C2(n220), .A(n1664), 
        .ZN(n1662) );
  AOI22_X1 U2114 ( .A1(n223), .A2(n4050), .B1(n29), .B2(n1200), .ZN(n1664) );
  OAI221_X1 U2115 ( .B1(n1665), .B2(n293), .C1(n945), .C2(n296), .A(n1666), 
        .ZN(n1661) );
  AOI22_X1 U2116 ( .A1(n299), .A2(n1302), .B1(n302), .B2(n4018), .ZN(n1666) );
  OAI211_X1 U2117 ( .C1(n529), .C2(n305), .A(n1667), .B(n1668), .ZN(n1660) );
  AOI221_X1 U2118 ( .B1(n307), .B2(n1161), .C1(n311), .C2(n4146), .A(n1669), 
        .ZN(n1668) );
  OAI22_X1 U2119 ( .A1(n625), .A2(n314), .B1(n1670), .B2(n317), .ZN(n1669) );
  AOI22_X1 U2120 ( .A1(n320), .A2(n4178), .B1(n323), .B2(n1059), .ZN(n1667) );
  NAND4_X1 U2121 ( .A1(n1674), .A2(n1671), .A3(n1673), .A4(n1672), .ZN(n1659)
         );
  AOI221_X1 U2122 ( .B1(n326), .B2(n4210), .C1(n329), .C2(n4242), .A(n1675), 
        .ZN(n1674) );
  OAI22_X1 U2123 ( .A1(n401), .A2(n333), .B1(n369), .B2(n20), .ZN(n1675) );
  AOI221_X1 U2124 ( .B1(n335), .B2(n4274), .C1(n338), .C2(n4306), .A(n1676), 
        .ZN(n1673) );
  OAI22_X1 U2125 ( .A1(n273), .A2(n342), .B1(n241), .B2(n344), .ZN(n1676) );
  AOI221_X1 U2126 ( .B1(n347), .B2(n782), .C1(n350), .C2(n816), .A(n1677), 
        .ZN(n1672) );
  OAI22_X1 U2127 ( .A1(n1678), .A2(n353), .B1(n1679), .B2(n356), .ZN(n1677) );
  OAI22_X1 U2128 ( .A1(n1681), .A2(n429), .B1(n1682), .B2(n5), .ZN(n1680) );
  OAI222_X1 U2129 ( .A1(n580), .A2(n208), .B1(n1683), .B2(n211), .C1(n3921), 
        .C2(n214), .ZN(n2556) );
  OAI221_X1 U2130 ( .B1(n850), .B2(n217), .C1(n1688), .C2(n220), .A(n1689), 
        .ZN(n1687) );
  AOI22_X1 U2131 ( .A1(n223), .A2(n4049), .B1(n225), .B2(n1201), .ZN(n1689) );
  OAI221_X1 U2132 ( .B1(n1690), .B2(n293), .C1(n946), .C2(n296), .A(n1691), 
        .ZN(n1686) );
  AOI22_X1 U2133 ( .A1(n299), .A2(n1303), .B1(n302), .B2(n4017), .ZN(n1691) );
  OAI211_X1 U2134 ( .C1(n530), .C2(n305), .A(n1692), .B(n1693), .ZN(n1685) );
  AOI221_X1 U2135 ( .B1(n308), .B2(n1162), .C1(n311), .C2(n4145), .A(n1694), 
        .ZN(n1693) );
  OAI22_X1 U2136 ( .A1(n626), .A2(n314), .B1(n1695), .B2(n317), .ZN(n1694) );
  AOI22_X1 U2137 ( .A1(n320), .A2(n4177), .B1(n323), .B2(n1060), .ZN(n1692) );
  NAND4_X1 U2138 ( .A1(n1696), .A2(n1697), .A3(n1698), .A4(n1699), .ZN(n1684)
         );
  AOI221_X1 U2139 ( .B1(n326), .B2(n4209), .C1(n329), .C2(n4241), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U2140 ( .A1(n402), .A2(n32), .B1(n370), .B2(n20), .ZN(n1700) );
  AOI221_X1 U2141 ( .B1(n335), .B2(n4273), .C1(n338), .C2(n4305), .A(n1701), 
        .ZN(n1698) );
  OAI22_X1 U2142 ( .A1(n274), .A2(n342), .B1(n242), .B2(n345), .ZN(n1701) );
  AOI221_X1 U2143 ( .B1(n347), .B2(n783), .C1(n350), .C2(n817), .A(n1702), 
        .ZN(n1697) );
  OAI22_X1 U2144 ( .A1(n1703), .A2(n353), .B1(n1704), .B2(n356), .ZN(n1702) );
  AOI221_X1 U2145 ( .B1(n422), .B2(n744), .C1(n426), .C2(n3953), .A(n1705), 
        .ZN(n1696) );
  OAI22_X1 U2146 ( .A1(n1706), .A2(n429), .B1(n1707), .B2(n23), .ZN(n1705) );
  OAI222_X1 U2147 ( .A1(n579), .A2(n208), .B1(n1708), .B2(n211), .C1(n3920), 
        .C2(n214), .ZN(n2555) );
  NOR4_X1 U2148 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .ZN(n1708)
         );
  OAI221_X1 U2149 ( .B1(n851), .B2(n217), .C1(n1713), .C2(n220), .A(n1714), 
        .ZN(n1712) );
  AOI22_X1 U2150 ( .A1(n223), .A2(n4048), .B1(n227), .B2(n1202), .ZN(n1714) );
  OAI221_X1 U2151 ( .B1(n1715), .B2(n293), .C1(n947), .C2(n296), .A(n1716), 
        .ZN(n1711) );
  AOI22_X1 U2152 ( .A1(n299), .A2(n1304), .B1(n302), .B2(n4016), .ZN(n1716) );
  OAI211_X1 U2153 ( .C1(n531), .C2(n305), .A(n1717), .B(n1718), .ZN(n1710) );
  AOI221_X1 U2154 ( .B1(n307), .B2(n1163), .C1(n311), .C2(n4144), .A(n1719), 
        .ZN(n1718) );
  OAI22_X1 U2155 ( .A1(n627), .A2(n314), .B1(n1720), .B2(n317), .ZN(n1719) );
  AOI22_X1 U2156 ( .A1(n320), .A2(n4176), .B1(n323), .B2(n1061), .ZN(n1717) );
  NAND4_X1 U2157 ( .A1(n1724), .A2(n1721), .A3(n1722), .A4(n1723), .ZN(n1709)
         );
  AOI221_X1 U2158 ( .B1(n326), .B2(n4208), .C1(n329), .C2(n4240), .A(n1725), 
        .ZN(n1724) );
  OAI22_X1 U2159 ( .A1(n403), .A2(n32), .B1(n371), .B2(n21), .ZN(n1725) );
  AOI221_X1 U2160 ( .B1(n335), .B2(n4272), .C1(n338), .C2(n4304), .A(n1726), 
        .ZN(n1723) );
  OAI22_X1 U2161 ( .A1(n275), .A2(n33), .B1(n243), .B2(n344), .ZN(n1726) );
  AOI221_X1 U2162 ( .B1(n347), .B2(n784), .C1(n350), .C2(n818), .A(n1727), 
        .ZN(n1722) );
  OAI22_X1 U2163 ( .A1(n1728), .A2(n353), .B1(n1729), .B2(n356), .ZN(n1727) );
  OAI22_X1 U2164 ( .A1(n1731), .A2(n429), .B1(n1732), .B2(n22), .ZN(n1730) );
  OAI222_X1 U2165 ( .A1(n578), .A2(n208), .B1(n1733), .B2(n211), .C1(n3919), 
        .C2(n214), .ZN(n2554) );
  OAI221_X1 U2166 ( .B1(n852), .B2(n217), .C1(n1738), .C2(n220), .A(n1739), 
        .ZN(n1737) );
  AOI22_X1 U2167 ( .A1(n223), .A2(n4047), .B1(n225), .B2(n1203), .ZN(n1739) );
  OAI221_X1 U2168 ( .B1(n1740), .B2(n293), .C1(n948), .C2(n296), .A(n1741), 
        .ZN(n1736) );
  AOI22_X1 U2169 ( .A1(n299), .A2(n1305), .B1(n302), .B2(n4015), .ZN(n1741) );
  OAI211_X1 U2170 ( .C1(n532), .C2(n305), .A(n1742), .B(n1743), .ZN(n1735) );
  AOI221_X1 U2171 ( .B1(n309), .B2(n1164), .C1(n311), .C2(n4143), .A(n1744), 
        .ZN(n1743) );
  OAI22_X1 U2172 ( .A1(n628), .A2(n314), .B1(n1745), .B2(n317), .ZN(n1744) );
  AOI22_X1 U2173 ( .A1(n320), .A2(n4175), .B1(n323), .B2(n1062), .ZN(n1742) );
  NAND4_X1 U2174 ( .A1(n1746), .A2(n1747), .A3(n1748), .A4(n1749), .ZN(n1734)
         );
  AOI221_X1 U2175 ( .B1(n326), .B2(n4207), .C1(n329), .C2(n4239), .A(n1750), 
        .ZN(n1749) );
  OAI22_X1 U2176 ( .A1(n404), .A2(n32), .B1(n372), .B2(n21), .ZN(n1750) );
  AOI221_X1 U2177 ( .B1(n335), .B2(n4271), .C1(n338), .C2(n4303), .A(n1751), 
        .ZN(n1748) );
  OAI22_X1 U2178 ( .A1(n276), .A2(n33), .B1(n244), .B2(n343), .ZN(n1751) );
  AOI221_X1 U2179 ( .B1(n347), .B2(n785), .C1(n350), .C2(n819), .A(n1752), 
        .ZN(n1747) );
  OAI22_X1 U2180 ( .A1(n1753), .A2(n353), .B1(n1754), .B2(n356), .ZN(n1752) );
  AOI221_X1 U2181 ( .B1(n423), .B2(n746), .C1(n426), .C2(n3951), .A(n1755), 
        .ZN(n1746) );
  OAI22_X1 U2182 ( .A1(n1756), .A2(n429), .B1(n1757), .B2(n23), .ZN(n1755) );
  OAI222_X1 U2183 ( .A1(n577), .A2(n208), .B1(n1758), .B2(n211), .C1(n3918), 
        .C2(n214), .ZN(n2553) );
  NOR4_X1 U2184 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(n1758)
         );
  OAI221_X1 U2185 ( .B1(n853), .B2(n217), .C1(n1763), .C2(n220), .A(n1764), 
        .ZN(n1762) );
  AOI22_X1 U2186 ( .A1(n223), .A2(n4046), .B1(n225), .B2(n1204), .ZN(n1764) );
  OAI221_X1 U2187 ( .B1(n1765), .B2(n293), .C1(n949), .C2(n296), .A(n1766), 
        .ZN(n1761) );
  AOI22_X1 U2188 ( .A1(n299), .A2(n1306), .B1(n302), .B2(n4014), .ZN(n1766) );
  OAI211_X1 U2189 ( .C1(n533), .C2(n305), .A(n1767), .B(n1768), .ZN(n1760) );
  AOI221_X1 U2190 ( .B1(n307), .B2(n1165), .C1(n311), .C2(n4142), .A(n1769), 
        .ZN(n1768) );
  OAI22_X1 U2191 ( .A1(n629), .A2(n314), .B1(n1770), .B2(n317), .ZN(n1769) );
  AOI22_X1 U2192 ( .A1(n320), .A2(n4174), .B1(n323), .B2(n1063), .ZN(n1767) );
  NAND4_X1 U2193 ( .A1(n1774), .A2(n1771), .A3(n1772), .A4(n1773), .ZN(n1759)
         );
  AOI221_X1 U2194 ( .B1(n326), .B2(n4206), .C1(n329), .C2(n4238), .A(n1775), 
        .ZN(n1774) );
  OAI22_X1 U2195 ( .A1(n405), .A2(n32), .B1(n373), .B2(n20), .ZN(n1775) );
  AOI221_X1 U2196 ( .B1(n335), .B2(n4270), .C1(n338), .C2(n4302), .A(n1776), 
        .ZN(n1773) );
  OAI22_X1 U2197 ( .A1(n277), .A2(n34), .B1(n245), .B2(n344), .ZN(n1776) );
  AOI221_X1 U2198 ( .B1(n347), .B2(n786), .C1(n350), .C2(n820), .A(n1777), 
        .ZN(n1772) );
  OAI22_X1 U2199 ( .A1(n1778), .A2(n353), .B1(n1779), .B2(n356), .ZN(n1777) );
  OAI22_X1 U2200 ( .A1(n1781), .A2(n429), .B1(n1782), .B2(n22), .ZN(n1780) );
  OAI222_X1 U2201 ( .A1(n576), .A2(n208), .B1(n1783), .B2(n211), .C1(n3917), 
        .C2(n214), .ZN(n2552) );
  OAI221_X1 U2202 ( .B1(n854), .B2(n217), .C1(n1788), .C2(n220), .A(n1789), 
        .ZN(n1787) );
  AOI22_X1 U2203 ( .A1(n223), .A2(n4045), .B1(n30), .B2(n1205), .ZN(n1789) );
  OAI221_X1 U2204 ( .B1(n1790), .B2(n293), .C1(n950), .C2(n296), .A(n1791), 
        .ZN(n1786) );
  AOI22_X1 U2205 ( .A1(n299), .A2(n1307), .B1(n302), .B2(n4013), .ZN(n1791) );
  OAI211_X1 U2206 ( .C1(n534), .C2(n305), .A(n1792), .B(n1793), .ZN(n1785) );
  AOI221_X1 U2207 ( .B1(n308), .B2(n1166), .C1(n311), .C2(n4141), .A(n1794), 
        .ZN(n1793) );
  OAI22_X1 U2208 ( .A1(n630), .A2(n314), .B1(n1795), .B2(n317), .ZN(n1794) );
  AOI22_X1 U2209 ( .A1(n320), .A2(n4173), .B1(n323), .B2(n1064), .ZN(n1792) );
  NAND4_X1 U2210 ( .A1(n1796), .A2(n1797), .A3(n1798), .A4(n1799), .ZN(n1784)
         );
  AOI221_X1 U2211 ( .B1(n326), .B2(n4205), .C1(n329), .C2(n4237), .A(n1800), 
        .ZN(n1799) );
  OAI22_X1 U2212 ( .A1(n406), .A2(n31), .B1(n374), .B2(n21), .ZN(n1800) );
  AOI221_X1 U2213 ( .B1(n335), .B2(n4269), .C1(n338), .C2(n4301), .A(n1801), 
        .ZN(n1798) );
  OAI22_X1 U2214 ( .A1(n278), .A2(n34), .B1(n246), .B2(n345), .ZN(n1801) );
  AOI221_X1 U2215 ( .B1(n347), .B2(n787), .C1(n350), .C2(n821), .A(n1802), 
        .ZN(n1797) );
  OAI22_X1 U2216 ( .A1(n1803), .A2(n353), .B1(n1804), .B2(n356), .ZN(n1802) );
  AOI221_X1 U2217 ( .B1(n422), .B2(n748), .C1(n426), .C2(n3949), .A(n1805), 
        .ZN(n1796) );
  OAI22_X1 U2218 ( .A1(n1806), .A2(n429), .B1(n1807), .B2(n22), .ZN(n1805) );
  OAI222_X1 U2219 ( .A1(n575), .A2(n208), .B1(n1808), .B2(n211), .C1(n3916), 
        .C2(n214), .ZN(n2551) );
  OAI221_X1 U2220 ( .B1(n855), .B2(n217), .C1(n1813), .C2(n220), .A(n1814), 
        .ZN(n1812) );
  AOI22_X1 U2221 ( .A1(n223), .A2(n4044), .B1(n226), .B2(n1206), .ZN(n1814) );
  OAI221_X1 U2222 ( .B1(n1815), .B2(n293), .C1(n951), .C2(n296), .A(n1816), 
        .ZN(n1811) );
  AOI22_X1 U2223 ( .A1(n299), .A2(n1308), .B1(n302), .B2(n4012), .ZN(n1816) );
  AOI221_X1 U2224 ( .B1(n309), .B2(n1167), .C1(n311), .C2(n4140), .A(n1819), 
        .ZN(n1818) );
  OAI22_X1 U2225 ( .A1(n631), .A2(n314), .B1(n1820), .B2(n317), .ZN(n1819) );
  AOI22_X1 U2226 ( .A1(n320), .A2(n4172), .B1(n323), .B2(n1065), .ZN(n1817) );
  NAND4_X1 U2227 ( .A1(n1824), .A2(n1821), .A3(n1822), .A4(n1823), .ZN(n1809)
         );
  AOI221_X1 U2228 ( .B1(n326), .B2(n4204), .C1(n329), .C2(n4236), .A(n1825), 
        .ZN(n1824) );
  OAI22_X1 U2229 ( .A1(n407), .A2(n332), .B1(n375), .B2(n20), .ZN(n1825) );
  AOI221_X1 U2230 ( .B1(n335), .B2(n4268), .C1(n338), .C2(n4300), .A(n1826), 
        .ZN(n1823) );
  OAI22_X1 U2231 ( .A1(n279), .A2(n341), .B1(n247), .B2(n344), .ZN(n1826) );
  AOI221_X1 U2232 ( .B1(n347), .B2(n788), .C1(n350), .C2(n822), .A(n1827), 
        .ZN(n1822) );
  OAI22_X1 U2233 ( .A1(n1828), .A2(n353), .B1(n1829), .B2(n356), .ZN(n1827) );
  OAI22_X1 U2234 ( .A1(n1831), .A2(n429), .B1(n1832), .B2(n22), .ZN(n1830) );
  OAI222_X1 U2235 ( .A1(n574), .A2(n208), .B1(n1833), .B2(n211), .C1(n3915), 
        .C2(n214), .ZN(n2550) );
  OAI221_X1 U2236 ( .B1(n856), .B2(n217), .C1(n1838), .C2(n220), .A(n1839), 
        .ZN(n1837) );
  AOI22_X1 U2237 ( .A1(n223), .A2(n4043), .B1(n29), .B2(n1207), .ZN(n1839) );
  OAI221_X1 U2238 ( .B1(n1840), .B2(n293), .C1(n952), .C2(n296), .A(n1841), 
        .ZN(n1836) );
  AOI22_X1 U2239 ( .A1(n299), .A2(n1309), .B1(n302), .B2(n4011), .ZN(n1841) );
  OAI211_X1 U2240 ( .C1(n536), .C2(n305), .A(n1842), .B(n1843), .ZN(n1835) );
  AOI221_X1 U2241 ( .B1(n309), .B2(n1168), .C1(n311), .C2(n4139), .A(n1844), 
        .ZN(n1843) );
  OAI22_X1 U2242 ( .A1(n632), .A2(n314), .B1(n1845), .B2(n317), .ZN(n1844) );
  AOI22_X1 U2243 ( .A1(n320), .A2(n4171), .B1(n323), .B2(n1066), .ZN(n1842) );
  NAND4_X1 U2244 ( .A1(n1846), .A2(n1847), .A3(n1848), .A4(n1849), .ZN(n1834)
         );
  AOI221_X1 U2245 ( .B1(n326), .B2(n4203), .C1(n329), .C2(n4235), .A(n1850), 
        .ZN(n1849) );
  OAI22_X1 U2246 ( .A1(n408), .A2(n31), .B1(n376), .B2(n21), .ZN(n1850) );
  AOI221_X1 U2247 ( .B1(n335), .B2(n4267), .C1(n338), .C2(n4299), .A(n1851), 
        .ZN(n1848) );
  OAI22_X1 U2248 ( .A1(n280), .A2(n341), .B1(n248), .B2(n343), .ZN(n1851) );
  AOI221_X1 U2249 ( .B1(n347), .B2(n789), .C1(n350), .C2(n823), .A(n1852), 
        .ZN(n1847) );
  OAI22_X1 U2250 ( .A1(n1853), .A2(n353), .B1(n1854), .B2(n356), .ZN(n1852) );
  AOI221_X1 U2251 ( .B1(n423), .B2(n750), .C1(n426), .C2(n3947), .A(n1855), 
        .ZN(n1846) );
  OAI22_X1 U2252 ( .A1(n1856), .A2(n429), .B1(n1857), .B2(n5), .ZN(n1855) );
  OAI222_X1 U2253 ( .A1(n573), .A2(n207), .B1(n1858), .B2(n210), .C1(n3914), 
        .C2(n214), .ZN(n2549) );
  NOR4_X1 U2254 ( .A1(n1859), .A2(n1860), .A3(n1861), .A4(n1862), .ZN(n1858)
         );
  OAI221_X1 U2255 ( .B1(n857), .B2(n216), .C1(n1863), .C2(n219), .A(n1864), 
        .ZN(n1862) );
  AOI22_X1 U2256 ( .A1(n222), .A2(n4042), .B1(n225), .B2(n1208), .ZN(n1864) );
  OAI221_X1 U2257 ( .B1(n1865), .B2(n228), .C1(n953), .C2(n295), .A(n1866), 
        .ZN(n1861) );
  AOI22_X1 U2258 ( .A1(n298), .A2(n1310), .B1(n301), .B2(n4010), .ZN(n1866) );
  OAI211_X1 U2259 ( .C1(n537), .C2(n304), .A(n1867), .B(n1868), .ZN(n1860) );
  AOI221_X1 U2260 ( .B1(n307), .B2(n1169), .C1(n310), .C2(n4138), .A(n1869), 
        .ZN(n1868) );
  OAI22_X1 U2261 ( .A1(n633), .A2(n313), .B1(n1870), .B2(n316), .ZN(n1869) );
  AOI22_X1 U2262 ( .A1(n319), .A2(n4170), .B1(n322), .B2(n1067), .ZN(n1867) );
  NAND4_X1 U2263 ( .A1(n1872), .A2(n1873), .A3(n1871), .A4(n1874), .ZN(n1859)
         );
  AOI221_X1 U2264 ( .B1(n325), .B2(n4202), .C1(n328), .C2(n4234), .A(n1875), 
        .ZN(n1874) );
  OAI22_X1 U2265 ( .A1(n409), .A2(n331), .B1(n377), .B2(n21), .ZN(n1875) );
  AOI221_X1 U2266 ( .B1(n334), .B2(n4266), .C1(n337), .C2(n4298), .A(n1876), 
        .ZN(n1873) );
  OAI22_X1 U2267 ( .A1(n281), .A2(n340), .B1(n249), .B2(n344), .ZN(n1876) );
  AOI221_X1 U2268 ( .B1(n346), .B2(n790), .C1(n349), .C2(n824), .A(n1877), 
        .ZN(n1872) );
  OAI22_X1 U2269 ( .A1(n1878), .A2(n352), .B1(n1879), .B2(n355), .ZN(n1877) );
  AOI221_X1 U2270 ( .B1(n424), .B2(n751), .C1(n425), .C2(n3946), .A(n1880), 
        .ZN(n1871) );
  OAI22_X1 U2271 ( .A1(n1881), .A2(n429), .B1(n1882), .B2(n5), .ZN(n1880) );
  OAI222_X1 U2272 ( .A1(n572), .A2(n207), .B1(n1883), .B2(n210), .C1(n3913), 
        .C2(n214), .ZN(n2548) );
  OAI221_X1 U2273 ( .B1(n858), .B2(n216), .C1(n1888), .C2(n219), .A(n1889), 
        .ZN(n1887) );
  AOI22_X1 U2274 ( .A1(n222), .A2(n4041), .B1(n225), .B2(n1209), .ZN(n1889) );
  OAI221_X1 U2275 ( .B1(n1890), .B2(n228), .C1(n954), .C2(n295), .A(n1891), 
        .ZN(n1886) );
  AOI22_X1 U2276 ( .A1(n298), .A2(n1311), .B1(n301), .B2(n4009), .ZN(n1891) );
  OAI211_X1 U2277 ( .C1(n538), .C2(n304), .A(n1892), .B(n1893), .ZN(n1885) );
  AOI221_X1 U2278 ( .B1(n308), .B2(n1170), .C1(n310), .C2(n4137), .A(n1894), 
        .ZN(n1893) );
  OAI22_X1 U2279 ( .A1(n634), .A2(n313), .B1(n1895), .B2(n316), .ZN(n1894) );
  AOI22_X1 U2280 ( .A1(n319), .A2(n4169), .B1(n322), .B2(n1068), .ZN(n1892) );
  NAND4_X1 U2281 ( .A1(n1896), .A2(n1897), .A3(n1898), .A4(n1899), .ZN(n1884)
         );
  AOI221_X1 U2282 ( .B1(n325), .B2(n4201), .C1(n328), .C2(n4233), .A(n1900), 
        .ZN(n1899) );
  OAI22_X1 U2283 ( .A1(n410), .A2(n32), .B1(n378), .B2(n20), .ZN(n1900) );
  AOI221_X1 U2284 ( .B1(n334), .B2(n4265), .C1(n337), .C2(n4297), .A(n1901), 
        .ZN(n1898) );
  OAI22_X1 U2285 ( .A1(n282), .A2(n340), .B1(n250), .B2(n345), .ZN(n1901) );
  AOI221_X1 U2286 ( .B1(n346), .B2(n791), .C1(n349), .C2(n825), .A(n1902), 
        .ZN(n1897) );
  OAI22_X1 U2287 ( .A1(n1903), .A2(n352), .B1(n1904), .B2(n355), .ZN(n1902) );
  AOI221_X1 U2288 ( .B1(n422), .B2(n752), .C1(n425), .C2(n3945), .A(n1905), 
        .ZN(n1896) );
  OAI22_X1 U2289 ( .A1(n1906), .A2(n428), .B1(n1907), .B2(n5), .ZN(n1905) );
  OAI222_X1 U2290 ( .A1(n571), .A2(n207), .B1(n1908), .B2(n210), .C1(n3912), 
        .C2(n213), .ZN(n2547) );
  NOR4_X1 U2291 ( .A1(n1909), .A2(n1910), .A3(n1911), .A4(n1912), .ZN(n1908)
         );
  OAI221_X1 U2292 ( .B1(n859), .B2(n216), .C1(n1913), .C2(n219), .A(n1914), 
        .ZN(n1912) );
  AOI22_X1 U2293 ( .A1(n222), .A2(n4040), .B1(n30), .B2(n1210), .ZN(n1914) );
  OAI221_X1 U2294 ( .B1(n1915), .B2(n228), .C1(n955), .C2(n295), .A(n1916), 
        .ZN(n1911) );
  AOI22_X1 U2295 ( .A1(n298), .A2(n1312), .B1(n301), .B2(n4008), .ZN(n1916) );
  OAI211_X1 U2296 ( .C1(n539), .C2(n304), .A(n1917), .B(n1918), .ZN(n1910) );
  AOI221_X1 U2297 ( .B1(n307), .B2(n1171), .C1(n310), .C2(n4136), .A(n1919), 
        .ZN(n1918) );
  OAI22_X1 U2298 ( .A1(n635), .A2(n313), .B1(n1920), .B2(n316), .ZN(n1919) );
  AOI22_X1 U2299 ( .A1(n319), .A2(n4168), .B1(n322), .B2(n1069), .ZN(n1917) );
  NAND4_X1 U2300 ( .A1(n1922), .A2(n1923), .A3(n1921), .A4(n1924), .ZN(n1909)
         );
  AOI221_X1 U2301 ( .B1(n325), .B2(n4200), .C1(n328), .C2(n4232), .A(n1925), 
        .ZN(n1924) );
  OAI22_X1 U2302 ( .A1(n411), .A2(n331), .B1(n379), .B2(n20), .ZN(n1925) );
  AOI221_X1 U2303 ( .B1(n334), .B2(n4264), .C1(n337), .C2(n4296), .A(n1926), 
        .ZN(n1923) );
  OAI22_X1 U2304 ( .A1(n283), .A2(n342), .B1(n251), .B2(n344), .ZN(n1926) );
  AOI221_X1 U2305 ( .B1(n346), .B2(n792), .C1(n349), .C2(n826), .A(n1927), 
        .ZN(n1922) );
  OAI22_X1 U2306 ( .A1(n1928), .A2(n352), .B1(n1929), .B2(n355), .ZN(n1927) );
  AOI221_X1 U2307 ( .B1(n424), .B2(n753), .C1(n425), .C2(n3944), .A(n1930), 
        .ZN(n1921) );
  OAI22_X1 U2308 ( .A1(n1931), .A2(n428), .B1(n1932), .B2(n23), .ZN(n1930) );
  OAI222_X1 U2309 ( .A1(n570), .A2(n207), .B1(n1933), .B2(n210), .C1(n3911), 
        .C2(n213), .ZN(n2546) );
  OAI221_X1 U2310 ( .B1(n860), .B2(n216), .C1(n1938), .C2(n219), .A(n1939), 
        .ZN(n1937) );
  AOI22_X1 U2311 ( .A1(n222), .A2(n4039), .B1(n30), .B2(n1211), .ZN(n1939) );
  OAI221_X1 U2312 ( .B1(n1940), .B2(n228), .C1(n956), .C2(n295), .A(n1941), 
        .ZN(n1936) );
  AOI22_X1 U2313 ( .A1(n298), .A2(n1313), .B1(n301), .B2(n4007), .ZN(n1941) );
  OAI211_X1 U2314 ( .C1(n540), .C2(n304), .A(n1942), .B(n1943), .ZN(n1935) );
  AOI221_X1 U2315 ( .B1(n309), .B2(n1172), .C1(n310), .C2(n4135), .A(n1944), 
        .ZN(n1943) );
  OAI22_X1 U2316 ( .A1(n636), .A2(n313), .B1(n1945), .B2(n316), .ZN(n1944) );
  AOI22_X1 U2317 ( .A1(n319), .A2(n4167), .B1(n322), .B2(n1070), .ZN(n1942) );
  NAND4_X1 U2318 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(n1934)
         );
  AOI221_X1 U2319 ( .B1(n325), .B2(n4199), .C1(n328), .C2(n4231), .A(n1950), 
        .ZN(n1949) );
  OAI22_X1 U2320 ( .A1(n412), .A2(n333), .B1(n380), .B2(n20), .ZN(n1950) );
  AOI221_X1 U2321 ( .B1(n334), .B2(n4263), .C1(n337), .C2(n4295), .A(n1951), 
        .ZN(n1948) );
  OAI22_X1 U2322 ( .A1(n284), .A2(n342), .B1(n252), .B2(n343), .ZN(n1951) );
  AOI221_X1 U2323 ( .B1(n346), .B2(n793), .C1(n349), .C2(n827), .A(n1952), 
        .ZN(n1947) );
  OAI22_X1 U2324 ( .A1(n1953), .A2(n352), .B1(n1954), .B2(n355), .ZN(n1952) );
  AOI221_X1 U2325 ( .B1(n423), .B2(n754), .C1(n425), .C2(n3943), .A(n1955), 
        .ZN(n1946) );
  OAI22_X1 U2326 ( .A1(n1956), .A2(n428), .B1(n1957), .B2(n23), .ZN(n1955) );
  OAI222_X1 U2327 ( .A1(n569), .A2(n207), .B1(n1958), .B2(n210), .C1(n3910), 
        .C2(n213), .ZN(n2545) );
  NOR4_X1 U2328 ( .A1(n1959), .A2(n1960), .A3(n1961), .A4(n1962), .ZN(n1958)
         );
  OAI221_X1 U2329 ( .B1(n861), .B2(n216), .C1(n1963), .C2(n219), .A(n1964), 
        .ZN(n1962) );
  AOI22_X1 U2330 ( .A1(n222), .A2(n4038), .B1(n29), .B2(n1212), .ZN(n1964) );
  OAI221_X1 U2331 ( .B1(n1965), .B2(n228), .C1(n957), .C2(n295), .A(n1966), 
        .ZN(n1961) );
  AOI22_X1 U2332 ( .A1(n298), .A2(n1314), .B1(n301), .B2(n4006), .ZN(n1966) );
  OAI211_X1 U2333 ( .C1(n541), .C2(n304), .A(n1967), .B(n1968), .ZN(n1960) );
  AOI221_X1 U2334 ( .B1(n307), .B2(n1173), .C1(n310), .C2(n4134), .A(n1969), 
        .ZN(n1968) );
  OAI22_X1 U2335 ( .A1(n637), .A2(n313), .B1(n1970), .B2(n316), .ZN(n1969) );
  AOI22_X1 U2336 ( .A1(n319), .A2(n4166), .B1(n322), .B2(n1071), .ZN(n1967) );
  NAND4_X1 U2337 ( .A1(n1972), .A2(n1973), .A3(n1971), .A4(n1974), .ZN(n1959)
         );
  AOI221_X1 U2338 ( .B1(n325), .B2(n4198), .C1(n328), .C2(n4230), .A(n1975), 
        .ZN(n1974) );
  OAI22_X1 U2339 ( .A1(n413), .A2(n331), .B1(n381), .B2(n21), .ZN(n1975) );
  AOI221_X1 U2340 ( .B1(n334), .B2(n4262), .C1(n337), .C2(n4294), .A(n1976), 
        .ZN(n1973) );
  OAI22_X1 U2341 ( .A1(n285), .A2(n33), .B1(n253), .B2(n344), .ZN(n1976) );
  AOI221_X1 U2342 ( .B1(n346), .B2(n794), .C1(n349), .C2(n828), .A(n1977), 
        .ZN(n1972) );
  OAI22_X1 U2343 ( .A1(n1978), .A2(n352), .B1(n1979), .B2(n355), .ZN(n1977) );
  AOI221_X1 U2344 ( .B1(n424), .B2(n755), .C1(n425), .C2(n3942), .A(n1980), 
        .ZN(n1971) );
  OAI22_X1 U2345 ( .A1(n1981), .A2(n428), .B1(n1982), .B2(n5), .ZN(n1980) );
  OAI222_X1 U2346 ( .A1(n568), .A2(n207), .B1(n1983), .B2(n210), .C1(n3909), 
        .C2(n213), .ZN(n2544) );
  OAI221_X1 U2347 ( .B1(n862), .B2(n216), .C1(n1988), .C2(n219), .A(n1989), 
        .ZN(n1987) );
  AOI22_X1 U2348 ( .A1(n222), .A2(n4037), .B1(n29), .B2(n1213), .ZN(n1989) );
  OAI221_X1 U2349 ( .B1(n1990), .B2(n228), .C1(n958), .C2(n295), .A(n1991), 
        .ZN(n1986) );
  AOI22_X1 U2350 ( .A1(n298), .A2(n1315), .B1(n301), .B2(n4005), .ZN(n1991) );
  OAI211_X1 U2351 ( .C1(n542), .C2(n304), .A(n1992), .B(n1993), .ZN(n1985) );
  AOI221_X1 U2352 ( .B1(n308), .B2(n1174), .C1(n310), .C2(n4133), .A(n1994), 
        .ZN(n1993) );
  OAI22_X1 U2353 ( .A1(n638), .A2(n313), .B1(n1995), .B2(n316), .ZN(n1994) );
  AOI22_X1 U2354 ( .A1(n319), .A2(n4165), .B1(n322), .B2(n1072), .ZN(n1992) );
  NAND4_X1 U2355 ( .A1(n1996), .A2(n1997), .A3(n1998), .A4(n1999), .ZN(n1984)
         );
  AOI221_X1 U2356 ( .B1(n325), .B2(n4197), .C1(n328), .C2(n4229), .A(n2000), 
        .ZN(n1999) );
  OAI22_X1 U2357 ( .A1(n414), .A2(n31), .B1(n382), .B2(n20), .ZN(n2000) );
  AOI221_X1 U2358 ( .B1(n334), .B2(n4261), .C1(n337), .C2(n4293), .A(n2001), 
        .ZN(n1998) );
  OAI22_X1 U2359 ( .A1(n286), .A2(n33), .B1(n254), .B2(n345), .ZN(n2001) );
  AOI221_X1 U2360 ( .B1(n346), .B2(n795), .C1(n349), .C2(n829), .A(n2002), 
        .ZN(n1997) );
  OAI22_X1 U2361 ( .A1(n2003), .A2(n352), .B1(n2004), .B2(n355), .ZN(n2002) );
  AOI221_X1 U2362 ( .B1(n422), .B2(n756), .C1(n425), .C2(n3941), .A(n2005), 
        .ZN(n1996) );
  OAI22_X1 U2363 ( .A1(n2006), .A2(n428), .B1(n2007), .B2(n23), .ZN(n2005) );
  OAI222_X1 U2364 ( .A1(n567), .A2(n207), .B1(n2008), .B2(n210), .C1(n3908), 
        .C2(n213), .ZN(n2543) );
  NOR4_X1 U2365 ( .A1(n2009), .A2(n2010), .A3(n2011), .A4(n2012), .ZN(n2008)
         );
  OAI221_X1 U2366 ( .B1(n863), .B2(n216), .C1(n2013), .C2(n219), .A(n2014), 
        .ZN(n2012) );
  AOI22_X1 U2367 ( .A1(n222), .A2(n4036), .B1(n227), .B2(n1214), .ZN(n2014) );
  OAI221_X1 U2368 ( .B1(n2015), .B2(n228), .C1(n959), .C2(n295), .A(n2016), 
        .ZN(n2011) );
  AOI22_X1 U2369 ( .A1(n298), .A2(n1316), .B1(n301), .B2(n4004), .ZN(n2016) );
  OAI211_X1 U2370 ( .C1(n543), .C2(n304), .A(n2017), .B(n2018), .ZN(n2010) );
  AOI221_X1 U2371 ( .B1(n307), .B2(n1175), .C1(n310), .C2(n4132), .A(n2019), 
        .ZN(n2018) );
  OAI22_X1 U2372 ( .A1(n639), .A2(n313), .B1(n2020), .B2(n316), .ZN(n2019) );
  AOI22_X1 U2373 ( .A1(n319), .A2(n4164), .B1(n322), .B2(n1073), .ZN(n2017) );
  NAND4_X1 U2374 ( .A1(n2022), .A2(n2023), .A3(n2021), .A4(n2024), .ZN(n2009)
         );
  AOI221_X1 U2375 ( .B1(n325), .B2(n4196), .C1(n328), .C2(n4228), .A(n2025), 
        .ZN(n2024) );
  OAI22_X1 U2376 ( .A1(n415), .A2(n331), .B1(n383), .B2(n20), .ZN(n2025) );
  AOI221_X1 U2377 ( .B1(n334), .B2(n4260), .C1(n337), .C2(n4292), .A(n2026), 
        .ZN(n2023) );
  OAI22_X1 U2378 ( .A1(n287), .A2(n34), .B1(n255), .B2(n344), .ZN(n2026) );
  AOI221_X1 U2379 ( .B1(n346), .B2(n796), .C1(n349), .C2(n830), .A(n2027), 
        .ZN(n2022) );
  OAI22_X1 U2380 ( .A1(n2028), .A2(n352), .B1(n2029), .B2(n355), .ZN(n2027) );
  AOI221_X1 U2381 ( .B1(n424), .B2(n757), .C1(n425), .C2(n3940), .A(n2030), 
        .ZN(n2021) );
  OAI22_X1 U2382 ( .A1(n2031), .A2(n428), .B1(n2032), .B2(n22), .ZN(n2030) );
  OAI222_X1 U2383 ( .A1(n566), .A2(n207), .B1(n2033), .B2(n210), .C1(n3907), 
        .C2(n213), .ZN(n2542) );
  OAI221_X1 U2384 ( .B1(n864), .B2(n216), .C1(n2038), .C2(n219), .A(n2039), 
        .ZN(n2037) );
  AOI22_X1 U2385 ( .A1(n222), .A2(n4035), .B1(n227), .B2(n1215), .ZN(n2039) );
  OAI221_X1 U2386 ( .B1(n2040), .B2(n228), .C1(n960), .C2(n295), .A(n2041), 
        .ZN(n2036) );
  AOI22_X1 U2387 ( .A1(n298), .A2(n1317), .B1(n301), .B2(n4003), .ZN(n2041) );
  OAI211_X1 U2388 ( .C1(n544), .C2(n304), .A(n2042), .B(n2043), .ZN(n2035) );
  AOI221_X1 U2389 ( .B1(n309), .B2(n1176), .C1(n310), .C2(n4131), .A(n2044), 
        .ZN(n2043) );
  OAI22_X1 U2390 ( .A1(n640), .A2(n313), .B1(n2045), .B2(n316), .ZN(n2044) );
  AOI22_X1 U2391 ( .A1(n319), .A2(n4163), .B1(n322), .B2(n1074), .ZN(n2042) );
  NAND4_X1 U2392 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .ZN(n2034)
         );
  AOI221_X1 U2393 ( .B1(n325), .B2(n4195), .C1(n328), .C2(n4227), .A(n2050), 
        .ZN(n2049) );
  OAI22_X1 U2394 ( .A1(n416), .A2(n332), .B1(n384), .B2(n21), .ZN(n2050) );
  AOI221_X1 U2395 ( .B1(n334), .B2(n4259), .C1(n337), .C2(n4291), .A(n2051), 
        .ZN(n2048) );
  OAI22_X1 U2396 ( .A1(n288), .A2(n34), .B1(n256), .B2(n343), .ZN(n2051) );
  AOI221_X1 U2397 ( .B1(n346), .B2(n797), .C1(n349), .C2(n831), .A(n2052), 
        .ZN(n2047) );
  OAI22_X1 U2398 ( .A1(n2053), .A2(n352), .B1(n2054), .B2(n355), .ZN(n2052) );
  AOI221_X1 U2399 ( .B1(n423), .B2(n758), .C1(n425), .C2(n3939), .A(n2055), 
        .ZN(n2046) );
  OAI22_X1 U2400 ( .A1(n2056), .A2(n428), .B1(n2057), .B2(n5), .ZN(n2055) );
  OAI222_X1 U2401 ( .A1(n565), .A2(n207), .B1(n2058), .B2(n210), .C1(n3906), 
        .C2(n213), .ZN(n2541) );
  OAI221_X1 U2402 ( .B1(n865), .B2(n216), .C1(n2063), .C2(n219), .A(n2064), 
        .ZN(n2062) );
  AOI22_X1 U2403 ( .A1(n222), .A2(n4034), .B1(n226), .B2(n1216), .ZN(n2064) );
  OAI221_X1 U2404 ( .B1(n2065), .B2(n228), .C1(n961), .C2(n295), .A(n2066), 
        .ZN(n2061) );
  AOI22_X1 U2405 ( .A1(n298), .A2(n1318), .B1(n301), .B2(n4002), .ZN(n2066) );
  OAI211_X1 U2406 ( .C1(n545), .C2(n304), .A(n2067), .B(n2068), .ZN(n2060) );
  AOI221_X1 U2407 ( .B1(n308), .B2(n1177), .C1(n310), .C2(n4130), .A(n2069), 
        .ZN(n2068) );
  OAI22_X1 U2408 ( .A1(n641), .A2(n313), .B1(n2070), .B2(n316), .ZN(n2069) );
  AOI22_X1 U2409 ( .A1(n319), .A2(n4162), .B1(n322), .B2(n1075), .ZN(n2067) );
  NAND4_X1 U2410 ( .A1(n2071), .A2(n2074), .A3(n2072), .A4(n2073), .ZN(n2059)
         );
  OAI22_X1 U2411 ( .A1(n417), .A2(n333), .B1(n385), .B2(n21), .ZN(n2075) );
  AOI221_X1 U2412 ( .B1(n334), .B2(n4258), .C1(n337), .C2(n4290), .A(n2076), 
        .ZN(n2073) );
  OAI22_X1 U2413 ( .A1(n289), .A2(n341), .B1(n257), .B2(n344), .ZN(n2076) );
  AOI221_X1 U2414 ( .B1(n346), .B2(n798), .C1(n349), .C2(n832), .A(n2077), 
        .ZN(n2072) );
  OAI22_X1 U2415 ( .A1(n2078), .A2(n352), .B1(n2079), .B2(n355), .ZN(n2077) );
  AOI221_X1 U2416 ( .B1(n422), .B2(n759), .C1(n425), .C2(n3938), .A(n2080), 
        .ZN(n2071) );
  OAI22_X1 U2417 ( .A1(n2081), .A2(n428), .B1(n2082), .B2(n5), .ZN(n2080) );
  OAI222_X1 U2418 ( .A1(n564), .A2(n207), .B1(n2083), .B2(n210), .C1(n3905), 
        .C2(n213), .ZN(n2540) );
  OAI221_X1 U2419 ( .B1(n866), .B2(n216), .C1(n2088), .C2(n219), .A(n2089), 
        .ZN(n2087) );
  AOI22_X1 U2420 ( .A1(n222), .A2(n4033), .B1(n227), .B2(n1217), .ZN(n2089) );
  OAI221_X1 U2421 ( .B1(n2090), .B2(n228), .C1(n962), .C2(n295), .A(n2091), 
        .ZN(n2086) );
  AOI22_X1 U2422 ( .A1(n298), .A2(n1319), .B1(n301), .B2(n4001), .ZN(n2091) );
  OAI211_X1 U2423 ( .C1(n546), .C2(n304), .A(n2092), .B(n2093), .ZN(n2085) );
  AOI221_X1 U2424 ( .B1(n308), .B2(n1178), .C1(n310), .C2(n4129), .A(n2094), 
        .ZN(n2093) );
  OAI22_X1 U2425 ( .A1(n642), .A2(n313), .B1(n2095), .B2(n316), .ZN(n2094) );
  AOI22_X1 U2426 ( .A1(n319), .A2(n4161), .B1(n322), .B2(n1076), .ZN(n2092) );
  NAND4_X1 U2427 ( .A1(n2096), .A2(n2097), .A3(n2098), .A4(n2099), .ZN(n2084)
         );
  AOI221_X1 U2428 ( .B1(n325), .B2(n4193), .C1(n328), .C2(n4225), .A(n2100), 
        .ZN(n2099) );
  OAI22_X1 U2429 ( .A1(n418), .A2(n31), .B1(n386), .B2(n21), .ZN(n2100) );
  AOI221_X1 U2430 ( .B1(n334), .B2(n4257), .C1(n337), .C2(n4289), .A(n2101), 
        .ZN(n2098) );
  OAI22_X1 U2431 ( .A1(n290), .A2(n341), .B1(n258), .B2(n343), .ZN(n2101) );
  OAI22_X1 U2432 ( .A1(n2103), .A2(n352), .B1(n2104), .B2(n355), .ZN(n2102) );
  AOI221_X1 U2433 ( .B1(n423), .B2(n760), .C1(n425), .C2(n3937), .A(n2105), 
        .ZN(n2096) );
  OAI22_X1 U2434 ( .A1(n2106), .A2(n428), .B1(n2107), .B2(n23), .ZN(n2105) );
  OAI222_X1 U2435 ( .A1(n563), .A2(n207), .B1(n2108), .B2(n210), .C1(n3904), 
        .C2(n213), .ZN(n2539) );
  OAI221_X1 U2436 ( .B1(n867), .B2(n216), .C1(n2113), .C2(n219), .A(n2114), 
        .ZN(n2112) );
  AOI22_X1 U2437 ( .A1(n222), .A2(n4032), .B1(n226), .B2(n1218), .ZN(n2114) );
  OAI221_X1 U2438 ( .B1(n2115), .B2(n228), .C1(n963), .C2(n295), .A(n2116), 
        .ZN(n2111) );
  AOI22_X1 U2439 ( .A1(n298), .A2(n1320), .B1(n301), .B2(n4000), .ZN(n2116) );
  AOI221_X1 U2440 ( .B1(n308), .B2(n1179), .C1(n310), .C2(n4128), .A(n2119), 
        .ZN(n2118) );
  OAI22_X1 U2441 ( .A1(n643), .A2(n313), .B1(n2120), .B2(n316), .ZN(n2119) );
  AOI22_X1 U2442 ( .A1(n319), .A2(n4160), .B1(n322), .B2(n1077), .ZN(n2117) );
  NAND4_X1 U2443 ( .A1(n2121), .A2(n2122), .A3(n2124), .A4(n2123), .ZN(n2109)
         );
  AOI221_X1 U2444 ( .B1(n325), .B2(n4192), .C1(n328), .C2(n4224), .A(n2125), 
        .ZN(n2124) );
  OAI22_X1 U2445 ( .A1(n419), .A2(n332), .B1(n387), .B2(n21), .ZN(n2125) );
  AOI221_X1 U2446 ( .B1(n334), .B2(n4256), .C1(n337), .C2(n4288), .A(n2126), 
        .ZN(n2123) );
  OAI22_X1 U2447 ( .A1(n291), .A2(n340), .B1(n259), .B2(n343), .ZN(n2126) );
  OAI22_X1 U2448 ( .A1(n2128), .A2(n352), .B1(n2129), .B2(n355), .ZN(n2127) );
  AOI221_X1 U2449 ( .B1(n422), .B2(n761), .C1(n425), .C2(n3936), .A(n2130), 
        .ZN(n2121) );
  OAI22_X1 U2450 ( .A1(n2131), .A2(n428), .B1(n2132), .B2(n22), .ZN(n2130) );
  OAI222_X1 U2451 ( .A1(n562), .A2(n207), .B1(n2133), .B2(n210), .C1(n3903), 
        .C2(n213), .ZN(n2538) );
  NAND2_X1 U2452 ( .A1(n213), .A2(n2134), .ZN(n1326) );
  OAI221_X1 U2453 ( .B1(n868), .B2(n216), .C1(n2139), .C2(n219), .A(n2140), 
        .ZN(n2138) );
  AOI22_X1 U2454 ( .A1(n222), .A2(n4031), .B1(n226), .B2(n1219), .ZN(n2140) );
  AND2_X1 U2455 ( .A1(n2141), .A2(n2142), .ZN(n1337) );
  AND2_X1 U2456 ( .A1(n2141), .A2(n2143), .ZN(n1336) );
  NAND2_X1 U2457 ( .A1(n2144), .A2(n2145), .ZN(n1334) );
  NAND2_X1 U2458 ( .A1(n2146), .A2(n2142), .ZN(n1332) );
  OAI221_X1 U2459 ( .B1(n2147), .B2(n228), .C1(n964), .C2(n295), .A(n2148), 
        .ZN(n2137) );
  AOI22_X1 U2460 ( .A1(n298), .A2(n1321), .B1(n301), .B2(n3999), .ZN(n2148) );
  AND2_X1 U2461 ( .A1(n2146), .A2(n2143), .ZN(n1343) );
  AND2_X1 U2462 ( .A1(n2146), .A2(n2145), .ZN(n1342) );
  NAND2_X1 U2463 ( .A1(n54), .A2(n2145), .ZN(n1340) );
  NAND2_X1 U2464 ( .A1(n54), .A2(n85), .ZN(n1339) );
  NOR3_X1 U2465 ( .A1(n2151), .A2(ADD_RS2[0]), .A3(n2150), .ZN(n2141) );
  OAI211_X1 U2466 ( .C1(n548), .C2(n304), .A(n2152), .B(n2153), .ZN(n2136) );
  AOI221_X1 U2467 ( .B1(n309), .B2(n1180), .C1(n310), .C2(n4127), .A(n2154), 
        .ZN(n2153) );
  OAI22_X1 U2468 ( .A1(n644), .A2(n313), .B1(n2155), .B2(n316), .ZN(n2154) );
  NAND2_X1 U2469 ( .A1(n2156), .A2(n2145), .ZN(n1352) );
  NAND2_X1 U2470 ( .A1(n2149), .A2(n2156), .ZN(n1350) );
  AND2_X1 U2471 ( .A1(n2144), .A2(n2142), .ZN(n1348) );
  AND2_X1 U2472 ( .A1(n2149), .A2(n2144), .ZN(n1347) );
  AOI22_X1 U2473 ( .A1(n319), .A2(n4159), .B1(n322), .B2(n1078), .ZN(n2152) );
  AND2_X1 U2474 ( .A1(n26), .A2(n18), .ZN(n1354) );
  AND2_X1 U2475 ( .A1(n26), .A2(n2142), .ZN(n1353) );
  NOR3_X1 U2476 ( .A1(ADD_RS2[0]), .A2(n86), .A3(ADD_RS2[3]), .ZN(n2156) );
  NAND2_X1 U2477 ( .A1(n2144), .A2(n18), .ZN(n1344) );
  NOR3_X1 U2478 ( .A1(n80), .A2(n2150), .A3(n77), .ZN(n2144) );
  NAND4_X1 U2479 ( .A1(n2157), .A2(n2158), .A3(n2160), .A4(n2159), .ZN(n2135)
         );
  AOI221_X1 U2480 ( .B1(n325), .B2(n4191), .C1(n328), .C2(n4223), .A(n2161), 
        .ZN(n2160) );
  OAI22_X1 U2481 ( .A1(n420), .A2(n333), .B1(n388), .B2(n20), .ZN(n2161) );
  NAND2_X1 U2482 ( .A1(n2162), .A2(n2149), .ZN(n1363) );
  NAND2_X1 U2483 ( .A1(n2163), .A2(n2149), .ZN(n1362) );
  AND2_X1 U2484 ( .A1(n19), .A2(n2145), .ZN(n1360) );
  AND2_X1 U2485 ( .A1(n2145), .A2(n35), .ZN(n1359) );
  AOI221_X1 U2486 ( .B1(n334), .B2(n4255), .C1(n337), .C2(n4287), .A(n2164), 
        .ZN(n2159) );
  OAI22_X1 U2487 ( .A1(n292), .A2(n340), .B1(n260), .B2(n345), .ZN(n2164) );
  NAND2_X1 U2488 ( .A1(n2162), .A2(n2143), .ZN(n1368) );
  NAND2_X1 U2489 ( .A1(n2163), .A2(n2143), .ZN(n1367) );
  AND2_X1 U2490 ( .A1(n2142), .A2(n19), .ZN(n1365) );
  NOR3_X1 U2491 ( .A1(n2151), .A2(ADD_RS2[4]), .A3(ADD_RS2[0]), .ZN(n2162) );
  AND2_X1 U2492 ( .A1(n2142), .A2(n35), .ZN(n1364) );
  NOR3_X1 U2493 ( .A1(n77), .A2(ADD_RS2[4]), .A3(n2151), .ZN(n2163) );
  OAI22_X1 U2494 ( .A1(n2166), .A2(n352), .B1(n2167), .B2(n355), .ZN(n2165) );
  NAND2_X1 U2495 ( .A1(n2168), .A2(n2145), .ZN(n1375) );
  NAND2_X1 U2496 ( .A1(n2169), .A2(n2145), .ZN(n1373) );
  AND2_X1 U2497 ( .A1(n79), .A2(n78), .ZN(n1370) );
  AND2_X1 U2498 ( .A1(n2169), .A2(n78), .ZN(n1369) );
  AOI221_X1 U2499 ( .B1(n422), .B2(n762), .C1(n425), .C2(n3935), .A(n2170), 
        .ZN(n2157) );
  OAI22_X1 U2500 ( .A1(n2171), .A2(n428), .B1(n2172), .B2(n22), .ZN(n2170) );
  NAND2_X1 U2501 ( .A1(n2168), .A2(n2142), .ZN(n1382) );
  NAND2_X1 U2502 ( .A1(n2169), .A2(n2142), .ZN(n1380) );
  NOR3_X1 U2503 ( .A1(ADD_RS2[0]), .A2(ADD_RS2[4]), .A3(ADD_RS2[3]), .ZN(n2169) );
  AND2_X1 U2504 ( .A1(n2146), .A2(n85), .ZN(n1377) );
  NOR2_X1 U2505 ( .A1(n2173), .A2(ADD_RS2[1]), .ZN(n2149) );
  INV_X1 U2506 ( .A(ADD_RS2[2]), .ZN(n2173) );
  NOR3_X1 U2507 ( .A1(n2150), .A2(n2151), .A3(n77), .ZN(n2146) );
  INV_X1 U2508 ( .A(ADD_RS2[3]), .ZN(n2151) );
  INV_X1 U2509 ( .A(ADD_RS2[4]), .ZN(n2150) );
  AND2_X1 U2510 ( .A1(n79), .A2(n2143), .ZN(n1376) );
  NOR2_X1 U2511 ( .A1(ADD_RS2[1]), .A2(ADD_RS2[2]), .ZN(n2143) );
  NAND2_X1 U2512 ( .A1(n2174), .A2(n213), .ZN(n1324) );
  AND3_X1 U2513 ( .A1(RD2), .A2(ENABLE), .A3(n715), .ZN(n1327) );
  INV_X1 U2514 ( .A(n2134), .ZN(n2174) );
  NAND4_X1 U2515 ( .A1(n2175), .A2(n2176), .A3(n2177), .A4(n2178), .ZN(n2134)
         );
  NOR3_X1 U2516 ( .A1(n2179), .A2(n1323), .A3(n2180), .ZN(n2178) );
  XNOR2_X1 U2517 ( .A(n1220), .B(n4), .ZN(n2180) );
  XNOR2_X1 U2518 ( .A(n1186), .B(n1), .ZN(n2179) );
  XNOR2_X1 U2519 ( .A(ADD_WR[3]), .B(n80), .ZN(n2177) );
  XNOR2_X1 U2520 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .ZN(n2176) );
  XNOR2_X1 U2521 ( .A(ADD_RS2[2]), .B(ADD_WR[2]), .ZN(n2175) );
  OAI222_X1 U2522 ( .A1(n593), .A2(n433), .B1(n2182), .B2(n436), .C1(n3902), 
        .C2(n439), .ZN(n2537) );
  NOR4_X1 U2523 ( .A1(n2185), .A2(n2186), .A3(n2187), .A4(n2188), .ZN(n2182)
         );
  OAI221_X1 U2524 ( .B1(n837), .B2(n442), .C1(n1333), .C2(n445), .A(n2191), 
        .ZN(n2188) );
  AOI22_X1 U2525 ( .A1(n448), .A2(n4062), .B1(n451), .B2(n1187), .ZN(n2191) );
  OAI221_X1 U2526 ( .B1(n1338), .B2(n454), .C1(n933), .C2(n457), .A(n2196), 
        .ZN(n2187) );
  AOI22_X1 U2527 ( .A1(n460), .A2(n1289), .B1(n463), .B2(n4030), .ZN(n2196) );
  OAI211_X1 U2528 ( .C1(n517), .C2(n466), .A(n2200), .B(n2201), .ZN(n2186) );
  AOI221_X1 U2529 ( .B1(n469), .B2(n1148), .C1(n472), .C2(n4158), .A(n2204), 
        .ZN(n2201) );
  OAI22_X1 U2530 ( .A1(n613), .A2(n475), .B1(n1351), .B2(n476), .ZN(n2204) );
  AOI22_X1 U2531 ( .A1(n481), .A2(n4190), .B1(n484), .B2(n1046), .ZN(n2200) );
  NAND4_X1 U2532 ( .A1(n2209), .A2(n2210), .A3(n2211), .A4(n2212), .ZN(n2185)
         );
  AOI221_X1 U2533 ( .B1(n487), .B2(n4222), .C1(n490), .C2(n4254), .A(n2215), 
        .ZN(n2212) );
  OAI22_X1 U2534 ( .A1(n389), .A2(n493), .B1(n357), .B2(n496), .ZN(n2215) );
  AOI221_X1 U2535 ( .B1(n499), .B2(n4286), .C1(n502), .C2(n4318), .A(n2220), 
        .ZN(n2211) );
  OAI22_X1 U2536 ( .A1(n261), .A2(n505), .B1(n229), .B2(n24), .ZN(n2220) );
  AOI221_X1 U2537 ( .B1(n508), .B2(n769), .C1(n511), .C2(n803), .A(n2225), 
        .ZN(n2210) );
  OAI22_X1 U2538 ( .A1(n1372), .A2(n514), .B1(n1374), .B2(n549), .ZN(n2225) );
  AOI221_X1 U2539 ( .B1(n552), .B2(n730), .C1(n555), .C2(n3966), .A(n2230), 
        .ZN(n2209) );
  OAI22_X1 U2540 ( .A1(n1379), .A2(n558), .B1(n1381), .B2(n561), .ZN(n2230) );
  OAI222_X1 U2541 ( .A1(n592), .A2(n433), .B1(n2233), .B2(n436), .C1(n3901), 
        .C2(n439), .ZN(n2536) );
  NOR4_X1 U2542 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2233)
         );
  OAI221_X1 U2543 ( .B1(n838), .B2(n442), .C1(n1388), .C2(n445), .A(n2238), 
        .ZN(n2237) );
  AOI22_X1 U2544 ( .A1(n448), .A2(n4061), .B1(n451), .B2(n1189), .ZN(n2238) );
  OAI221_X1 U2545 ( .B1(n1390), .B2(n454), .C1(n934), .C2(n457), .A(n2239), 
        .ZN(n2236) );
  AOI22_X1 U2546 ( .A1(n460), .A2(n1291), .B1(n463), .B2(n4029), .ZN(n2239) );
  OAI211_X1 U2547 ( .C1(n518), .C2(n466), .A(n2240), .B(n2241), .ZN(n2235) );
  AOI221_X1 U2548 ( .B1(n469), .B2(n1150), .C1(n472), .C2(n4157), .A(n2242), 
        .ZN(n2241) );
  OAI22_X1 U2549 ( .A1(n614), .A2(n473), .B1(n1395), .B2(n477), .ZN(n2242) );
  AOI22_X1 U2550 ( .A1(n481), .A2(n4189), .B1(n484), .B2(n1048), .ZN(n2240) );
  NAND4_X1 U2551 ( .A1(n2243), .A2(n2244), .A3(n2245), .A4(n2246), .ZN(n2234)
         );
  AOI221_X1 U2552 ( .B1(n487), .B2(n4221), .C1(n490), .C2(n4253), .A(n2247), 
        .ZN(n2246) );
  OAI22_X1 U2553 ( .A1(n390), .A2(n493), .B1(n358), .B2(n496), .ZN(n2247) );
  AOI221_X1 U2554 ( .B1(n499), .B2(n4285), .C1(n502), .C2(n4317), .A(n2248), 
        .ZN(n2245) );
  OAI22_X1 U2555 ( .A1(n262), .A2(n505), .B1(n230), .B2(n25), .ZN(n2248) );
  AOI221_X1 U2556 ( .B1(n508), .B2(n771), .C1(n511), .C2(n805), .A(n2249), 
        .ZN(n2244) );
  OAI22_X1 U2557 ( .A1(n1403), .A2(n514), .B1(n1404), .B2(n549), .ZN(n2249) );
  AOI221_X1 U2558 ( .B1(n552), .B2(n732), .C1(n555), .C2(n3965), .A(n2250), 
        .ZN(n2243) );
  OAI22_X1 U2559 ( .A1(n1406), .A2(n558), .B1(n1407), .B2(n561), .ZN(n2250) );
  OAI222_X1 U2560 ( .A1(n591), .A2(n433), .B1(n2251), .B2(n436), .C1(n3900), 
        .C2(n439), .ZN(n2535) );
  NOR4_X1 U2561 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  OAI221_X1 U2562 ( .B1(n839), .B2(n442), .C1(n1413), .C2(n445), .A(n2256), 
        .ZN(n2255) );
  AOI22_X1 U2563 ( .A1(n448), .A2(n4060), .B1(n451), .B2(n1190), .ZN(n2256) );
  OAI221_X1 U2564 ( .B1(n1415), .B2(n454), .C1(n935), .C2(n457), .A(n2257), 
        .ZN(n2254) );
  AOI22_X1 U2565 ( .A1(n460), .A2(n1292), .B1(n463), .B2(n4028), .ZN(n2257) );
  OAI211_X1 U2566 ( .C1(n519), .C2(n466), .A(n2258), .B(n2259), .ZN(n2253) );
  AOI221_X1 U2567 ( .B1(n469), .B2(n1151), .C1(n472), .C2(n4156), .A(n2260), 
        .ZN(n2259) );
  OAI22_X1 U2568 ( .A1(n615), .A2(n28), .B1(n1420), .B2(n478), .ZN(n2260) );
  AOI22_X1 U2569 ( .A1(n481), .A2(n4188), .B1(n484), .B2(n1049), .ZN(n2258) );
  NAND4_X1 U2570 ( .A1(n2261), .A2(n2262), .A3(n2263), .A4(n2264), .ZN(n2252)
         );
  AOI221_X1 U2571 ( .B1(n487), .B2(n4220), .C1(n490), .C2(n4252), .A(n2265), 
        .ZN(n2264) );
  OAI22_X1 U2572 ( .A1(n391), .A2(n493), .B1(n359), .B2(n496), .ZN(n2265) );
  AOI221_X1 U2573 ( .B1(n499), .B2(n4284), .C1(n502), .C2(n4316), .A(n2266), 
        .ZN(n2263) );
  OAI22_X1 U2574 ( .A1(n263), .A2(n505), .B1(n231), .B2(n24), .ZN(n2266) );
  AOI221_X1 U2575 ( .B1(n508), .B2(n772), .C1(n511), .C2(n806), .A(n2267), 
        .ZN(n2262) );
  OAI22_X1 U2576 ( .A1(n1428), .A2(n514), .B1(n1429), .B2(n549), .ZN(n2267) );
  AOI221_X1 U2577 ( .B1(n552), .B2(n733), .C1(n555), .C2(n3964), .A(n2268), 
        .ZN(n2261) );
  OAI22_X1 U2578 ( .A1(n1431), .A2(n558), .B1(n1432), .B2(n561), .ZN(n2268) );
  OAI222_X1 U2579 ( .A1(n590), .A2(n433), .B1(n2269), .B2(n436), .C1(n3899), 
        .C2(n439), .ZN(n2534) );
  NOR4_X1 U2580 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n2269)
         );
  OAI221_X1 U2581 ( .B1(n840), .B2(n442), .C1(n1438), .C2(n445), .A(n2274), 
        .ZN(n2273) );
  AOI22_X1 U2582 ( .A1(n448), .A2(n4059), .B1(n451), .B2(n1191), .ZN(n2274) );
  OAI221_X1 U2583 ( .B1(n1440), .B2(n454), .C1(n936), .C2(n457), .A(n2275), 
        .ZN(n2272) );
  AOI22_X1 U2584 ( .A1(n460), .A2(n1293), .B1(n463), .B2(n4027), .ZN(n2275) );
  OAI211_X1 U2585 ( .C1(n520), .C2(n466), .A(n2276), .B(n2277), .ZN(n2271) );
  AOI221_X1 U2586 ( .B1(n469), .B2(n1152), .C1(n472), .C2(n4155), .A(n2278), 
        .ZN(n2277) );
  OAI22_X1 U2587 ( .A1(n616), .A2(n27), .B1(n1445), .B2(n476), .ZN(n2278) );
  AOI22_X1 U2588 ( .A1(n481), .A2(n4187), .B1(n484), .B2(n1050), .ZN(n2276) );
  NAND4_X1 U2589 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2270)
         );
  AOI221_X1 U2590 ( .B1(n487), .B2(n4219), .C1(n490), .C2(n4251), .A(n2283), 
        .ZN(n2282) );
  OAI22_X1 U2591 ( .A1(n392), .A2(n493), .B1(n360), .B2(n496), .ZN(n2283) );
  AOI221_X1 U2592 ( .B1(n499), .B2(n4283), .C1(n502), .C2(n4315), .A(n2284), 
        .ZN(n2281) );
  OAI22_X1 U2593 ( .A1(n264), .A2(n505), .B1(n232), .B2(n25), .ZN(n2284) );
  AOI221_X1 U2594 ( .B1(n508), .B2(n773), .C1(n511), .C2(n807), .A(n2285), 
        .ZN(n2280) );
  OAI22_X1 U2595 ( .A1(n1453), .A2(n514), .B1(n1454), .B2(n549), .ZN(n2285) );
  AOI221_X1 U2596 ( .B1(n552), .B2(n734), .C1(n555), .C2(n3963), .A(n2286), 
        .ZN(n2279) );
  OAI22_X1 U2597 ( .A1(n1456), .A2(n558), .B1(n1457), .B2(n561), .ZN(n2286) );
  OAI222_X1 U2598 ( .A1(n589), .A2(n433), .B1(n2287), .B2(n436), .C1(n3898), 
        .C2(n439), .ZN(n2533) );
  NOR4_X1 U2599 ( .A1(n2288), .A2(n2289), .A3(n2290), .A4(n2291), .ZN(n2287)
         );
  OAI221_X1 U2600 ( .B1(n841), .B2(n442), .C1(n1463), .C2(n445), .A(n2292), 
        .ZN(n2291) );
  AOI22_X1 U2601 ( .A1(n448), .A2(n4058), .B1(n451), .B2(n1192), .ZN(n2292) );
  OAI221_X1 U2602 ( .B1(n1465), .B2(n454), .C1(n937), .C2(n457), .A(n2293), 
        .ZN(n2290) );
  AOI22_X1 U2603 ( .A1(n460), .A2(n1294), .B1(n463), .B2(n4026), .ZN(n2293) );
  OAI211_X1 U2604 ( .C1(n521), .C2(n466), .A(n2294), .B(n2295), .ZN(n2289) );
  AOI221_X1 U2605 ( .B1(n469), .B2(n1153), .C1(n472), .C2(n4154), .A(n2296), 
        .ZN(n2295) );
  OAI22_X1 U2606 ( .A1(n617), .A2(n475), .B1(n1470), .B2(n478), .ZN(n2296) );
  AOI22_X1 U2607 ( .A1(n481), .A2(n4186), .B1(n484), .B2(n1051), .ZN(n2294) );
  NAND4_X1 U2608 ( .A1(n2297), .A2(n2298), .A3(n2299), .A4(n2300), .ZN(n2288)
         );
  AOI221_X1 U2609 ( .B1(n487), .B2(n4218), .C1(n490), .C2(n4250), .A(n2301), 
        .ZN(n2300) );
  OAI22_X1 U2610 ( .A1(n393), .A2(n493), .B1(n361), .B2(n496), .ZN(n2301) );
  AOI221_X1 U2611 ( .B1(n499), .B2(n4282), .C1(n502), .C2(n4314), .A(n2302), 
        .ZN(n2299) );
  OAI22_X1 U2612 ( .A1(n265), .A2(n505), .B1(n233), .B2(n24), .ZN(n2302) );
  AOI221_X1 U2613 ( .B1(n508), .B2(n774), .C1(n511), .C2(n808), .A(n2303), 
        .ZN(n2298) );
  OAI22_X1 U2614 ( .A1(n1478), .A2(n514), .B1(n1479), .B2(n549), .ZN(n2303) );
  AOI221_X1 U2615 ( .B1(n552), .B2(n735), .C1(n555), .C2(n3962), .A(n2304), 
        .ZN(n2297) );
  OAI22_X1 U2616 ( .A1(n1481), .A2(n558), .B1(n1482), .B2(n561), .ZN(n2304) );
  OAI222_X1 U2617 ( .A1(n588), .A2(n433), .B1(n2305), .B2(n436), .C1(n3897), 
        .C2(n439), .ZN(n2532) );
  NOR4_X1 U2618 ( .A1(n2306), .A2(n2307), .A3(n2308), .A4(n2309), .ZN(n2305)
         );
  OAI221_X1 U2619 ( .B1(n842), .B2(n442), .C1(n1488), .C2(n445), .A(n2310), 
        .ZN(n2309) );
  AOI22_X1 U2620 ( .A1(n448), .A2(n4057), .B1(n451), .B2(n1193), .ZN(n2310) );
  OAI221_X1 U2621 ( .B1(n1490), .B2(n454), .C1(n938), .C2(n457), .A(n2311), 
        .ZN(n2308) );
  AOI22_X1 U2622 ( .A1(n460), .A2(n1295), .B1(n463), .B2(n4025), .ZN(n2311) );
  OAI211_X1 U2623 ( .C1(n522), .C2(n466), .A(n2312), .B(n2313), .ZN(n2307) );
  AOI221_X1 U2624 ( .B1(n469), .B2(n1154), .C1(n472), .C2(n4153), .A(n2314), 
        .ZN(n2313) );
  OAI22_X1 U2625 ( .A1(n618), .A2(n473), .B1(n1495), .B2(n478), .ZN(n2314) );
  AOI22_X1 U2626 ( .A1(n481), .A2(n4185), .B1(n484), .B2(n1052), .ZN(n2312) );
  NAND4_X1 U2627 ( .A1(n2315), .A2(n2316), .A3(n2317), .A4(n2318), .ZN(n2306)
         );
  AOI221_X1 U2628 ( .B1(n487), .B2(n4217), .C1(n490), .C2(n4249), .A(n2319), 
        .ZN(n2318) );
  OAI22_X1 U2629 ( .A1(n394), .A2(n493), .B1(n362), .B2(n496), .ZN(n2319) );
  AOI221_X1 U2630 ( .B1(n499), .B2(n4281), .C1(n502), .C2(n4313), .A(n2320), 
        .ZN(n2317) );
  OAI22_X1 U2631 ( .A1(n266), .A2(n505), .B1(n234), .B2(n25), .ZN(n2320) );
  AOI221_X1 U2632 ( .B1(n508), .B2(n775), .C1(n511), .C2(n809), .A(n2321), 
        .ZN(n2316) );
  OAI22_X1 U2633 ( .A1(n1503), .A2(n514), .B1(n1504), .B2(n549), .ZN(n2321) );
  AOI221_X1 U2634 ( .B1(n552), .B2(n736), .C1(n555), .C2(n3961), .A(n2322), 
        .ZN(n2315) );
  OAI22_X1 U2635 ( .A1(n1506), .A2(n558), .B1(n1507), .B2(n561), .ZN(n2322) );
  OAI222_X1 U2636 ( .A1(n587), .A2(n433), .B1(n2323), .B2(n436), .C1(n3896), 
        .C2(n439), .ZN(n2531) );
  NOR4_X1 U2637 ( .A1(n2324), .A2(n2325), .A3(n2326), .A4(n2327), .ZN(n2323)
         );
  OAI221_X1 U2638 ( .B1(n843), .B2(n442), .C1(n1513), .C2(n445), .A(n2328), 
        .ZN(n2327) );
  AOI22_X1 U2639 ( .A1(n448), .A2(n4056), .B1(n451), .B2(n1194), .ZN(n2328) );
  OAI221_X1 U2640 ( .B1(n1515), .B2(n454), .C1(n939), .C2(n457), .A(n2329), 
        .ZN(n2326) );
  AOI22_X1 U2641 ( .A1(n460), .A2(n1296), .B1(n463), .B2(n4024), .ZN(n2329) );
  OAI211_X1 U2642 ( .C1(n523), .C2(n466), .A(n2330), .B(n2331), .ZN(n2325) );
  AOI221_X1 U2643 ( .B1(n469), .B2(n1155), .C1(n472), .C2(n4152), .A(n2332), 
        .ZN(n2331) );
  OAI22_X1 U2644 ( .A1(n619), .A2(n28), .B1(n1520), .B2(n476), .ZN(n2332) );
  AOI22_X1 U2645 ( .A1(n481), .A2(n4184), .B1(n484), .B2(n1053), .ZN(n2330) );
  NAND4_X1 U2646 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(n2324)
         );
  AOI221_X1 U2647 ( .B1(n487), .B2(n4216), .C1(n490), .C2(n4248), .A(n2337), 
        .ZN(n2336) );
  OAI22_X1 U2648 ( .A1(n395), .A2(n493), .B1(n363), .B2(n496), .ZN(n2337) );
  AOI221_X1 U2649 ( .B1(n499), .B2(n4280), .C1(n502), .C2(n4312), .A(n2338), 
        .ZN(n2335) );
  OAI22_X1 U2650 ( .A1(n267), .A2(n505), .B1(n235), .B2(n24), .ZN(n2338) );
  AOI221_X1 U2651 ( .B1(n508), .B2(n776), .C1(n511), .C2(n810), .A(n2339), 
        .ZN(n2334) );
  OAI22_X1 U2652 ( .A1(n1528), .A2(n514), .B1(n1529), .B2(n549), .ZN(n2339) );
  AOI221_X1 U2653 ( .B1(n552), .B2(n737), .C1(n555), .C2(n3960), .A(n2340), 
        .ZN(n2333) );
  OAI22_X1 U2654 ( .A1(n1531), .A2(n558), .B1(n1532), .B2(n561), .ZN(n2340) );
  OAI222_X1 U2655 ( .A1(n586), .A2(n433), .B1(n2341), .B2(n436), .C1(n3895), 
        .C2(n439), .ZN(n2530) );
  NOR4_X1 U2656 ( .A1(n2342), .A2(n2343), .A3(n2344), .A4(n2345), .ZN(n2341)
         );
  OAI221_X1 U2657 ( .B1(n844), .B2(n442), .C1(n1538), .C2(n445), .A(n2346), 
        .ZN(n2345) );
  AOI22_X1 U2658 ( .A1(n448), .A2(n4055), .B1(n451), .B2(n1195), .ZN(n2346) );
  OAI221_X1 U2659 ( .B1(n1540), .B2(n454), .C1(n940), .C2(n457), .A(n2347), 
        .ZN(n2344) );
  AOI22_X1 U2660 ( .A1(n460), .A2(n1297), .B1(n463), .B2(n4023), .ZN(n2347) );
  OAI211_X1 U2661 ( .C1(n524), .C2(n466), .A(n2348), .B(n2349), .ZN(n2343) );
  AOI221_X1 U2662 ( .B1(n469), .B2(n1156), .C1(n472), .C2(n4151), .A(n2350), 
        .ZN(n2349) );
  OAI22_X1 U2663 ( .A1(n620), .A2(n27), .B1(n1545), .B2(n478), .ZN(n2350) );
  AOI22_X1 U2664 ( .A1(n481), .A2(n4183), .B1(n484), .B2(n1054), .ZN(n2348) );
  NAND4_X1 U2665 ( .A1(n2351), .A2(n2352), .A3(n2353), .A4(n2354), .ZN(n2342)
         );
  AOI221_X1 U2666 ( .B1(n487), .B2(n4215), .C1(n490), .C2(n4247), .A(n2355), 
        .ZN(n2354) );
  OAI22_X1 U2667 ( .A1(n396), .A2(n493), .B1(n364), .B2(n496), .ZN(n2355) );
  AOI221_X1 U2668 ( .B1(n499), .B2(n4279), .C1(n502), .C2(n4311), .A(n2356), 
        .ZN(n2353) );
  OAI22_X1 U2669 ( .A1(n268), .A2(n505), .B1(n236), .B2(n25), .ZN(n2356) );
  AOI221_X1 U2670 ( .B1(n508), .B2(n777), .C1(n511), .C2(n811), .A(n2357), 
        .ZN(n2352) );
  OAI22_X1 U2671 ( .A1(n1553), .A2(n514), .B1(n1554), .B2(n549), .ZN(n2357) );
  AOI221_X1 U2672 ( .B1(n552), .B2(n738), .C1(n555), .C2(n3959), .A(n2358), 
        .ZN(n2351) );
  OAI22_X1 U2673 ( .A1(n1556), .A2(n558), .B1(n1557), .B2(n561), .ZN(n2358) );
  OAI222_X1 U2674 ( .A1(n585), .A2(n432), .B1(n2359), .B2(n435), .C1(n3894), 
        .C2(n439), .ZN(n2529) );
  NOR4_X1 U2675 ( .A1(n2360), .A2(n2361), .A3(n2362), .A4(n2363), .ZN(n2359)
         );
  OAI221_X1 U2676 ( .B1(n845), .B2(n441), .C1(n1563), .C2(n444), .A(n2364), 
        .ZN(n2363) );
  AOI22_X1 U2677 ( .A1(n447), .A2(n4054), .B1(n450), .B2(n1196), .ZN(n2364) );
  OAI221_X1 U2678 ( .B1(n1565), .B2(n453), .C1(n941), .C2(n456), .A(n2365), 
        .ZN(n2362) );
  AOI22_X1 U2679 ( .A1(n459), .A2(n1298), .B1(n462), .B2(n4022), .ZN(n2365) );
  OAI211_X1 U2680 ( .C1(n525), .C2(n465), .A(n2366), .B(n2367), .ZN(n2361) );
  AOI221_X1 U2681 ( .B1(n468), .B2(n1157), .C1(n471), .C2(n4150), .A(n2368), 
        .ZN(n2367) );
  OAI22_X1 U2682 ( .A1(n621), .A2(n474), .B1(n1570), .B2(n477), .ZN(n2368) );
  AOI22_X1 U2683 ( .A1(n480), .A2(n4182), .B1(n483), .B2(n1055), .ZN(n2366) );
  NAND4_X1 U2684 ( .A1(n2369), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n2360)
         );
  AOI221_X1 U2685 ( .B1(n486), .B2(n4214), .C1(n489), .C2(n4246), .A(n2373), 
        .ZN(n2372) );
  OAI22_X1 U2686 ( .A1(n397), .A2(n492), .B1(n365), .B2(n496), .ZN(n2373) );
  AOI221_X1 U2687 ( .B1(n498), .B2(n4278), .C1(n501), .C2(n4310), .A(n2374), 
        .ZN(n2371) );
  OAI22_X1 U2688 ( .A1(n269), .A2(n504), .B1(n237), .B2(n25), .ZN(n2374) );
  AOI221_X1 U2689 ( .B1(n507), .B2(n778), .C1(n510), .C2(n812), .A(n2375), 
        .ZN(n2370) );
  OAI22_X1 U2690 ( .A1(n1578), .A2(n513), .B1(n1579), .B2(n549), .ZN(n2375) );
  AOI221_X1 U2691 ( .B1(n551), .B2(n739), .C1(n554), .C2(n3958), .A(n2376), 
        .ZN(n2369) );
  OAI22_X1 U2692 ( .A1(n1581), .A2(n557), .B1(n1582), .B2(n560), .ZN(n2376) );
  OAI222_X1 U2693 ( .A1(n584), .A2(n432), .B1(n2377), .B2(n435), .C1(n3893), 
        .C2(n439), .ZN(n2528) );
  NOR4_X1 U2694 ( .A1(n2378), .A2(n2379), .A3(n2380), .A4(n2381), .ZN(n2377)
         );
  OAI221_X1 U2695 ( .B1(n846), .B2(n441), .C1(n1588), .C2(n444), .A(n2382), 
        .ZN(n2381) );
  AOI22_X1 U2696 ( .A1(n447), .A2(n4053), .B1(n450), .B2(n1197), .ZN(n2382) );
  OAI221_X1 U2697 ( .B1(n1590), .B2(n453), .C1(n942), .C2(n456), .A(n2383), 
        .ZN(n2380) );
  AOI22_X1 U2698 ( .A1(n459), .A2(n1299), .B1(n462), .B2(n4021), .ZN(n2383) );
  OAI211_X1 U2699 ( .C1(n526), .C2(n465), .A(n2384), .B(n2385), .ZN(n2379) );
  AOI221_X1 U2700 ( .B1(n468), .B2(n1158), .C1(n471), .C2(n4149), .A(n2386), 
        .ZN(n2385) );
  OAI22_X1 U2701 ( .A1(n622), .A2(n474), .B1(n1595), .B2(n477), .ZN(n2386) );
  AOI22_X1 U2702 ( .A1(n480), .A2(n4181), .B1(n483), .B2(n1056), .ZN(n2384) );
  NAND4_X1 U2703 ( .A1(n2387), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n2378)
         );
  AOI221_X1 U2704 ( .B1(n486), .B2(n4213), .C1(n489), .C2(n4245), .A(n2391), 
        .ZN(n2390) );
  OAI22_X1 U2705 ( .A1(n398), .A2(n492), .B1(n366), .B2(n495), .ZN(n2391) );
  AOI221_X1 U2706 ( .B1(n498), .B2(n4277), .C1(n501), .C2(n4309), .A(n2392), 
        .ZN(n2389) );
  OAI22_X1 U2707 ( .A1(n270), .A2(n504), .B1(n238), .B2(n24), .ZN(n2392) );
  AOI221_X1 U2708 ( .B1(n507), .B2(n779), .C1(n510), .C2(n813), .A(n2393), 
        .ZN(n2388) );
  OAI22_X1 U2709 ( .A1(n1603), .A2(n513), .B1(n1604), .B2(n516), .ZN(n2393) );
  AOI221_X1 U2710 ( .B1(n551), .B2(n740), .C1(n554), .C2(n3957), .A(n2394), 
        .ZN(n2387) );
  OAI22_X1 U2711 ( .A1(n1606), .A2(n557), .B1(n1607), .B2(n560), .ZN(n2394) );
  OAI222_X1 U2712 ( .A1(n583), .A2(n432), .B1(n2395), .B2(n435), .C1(n3892), 
        .C2(n438), .ZN(n2527) );
  NOR4_X1 U2713 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(n2395)
         );
  OAI221_X1 U2714 ( .B1(n847), .B2(n441), .C1(n1613), .C2(n444), .A(n2400), 
        .ZN(n2399) );
  AOI22_X1 U2715 ( .A1(n447), .A2(n4052), .B1(n450), .B2(n1198), .ZN(n2400) );
  OAI221_X1 U2716 ( .B1(n1615), .B2(n453), .C1(n943), .C2(n456), .A(n2401), 
        .ZN(n2398) );
  AOI22_X1 U2717 ( .A1(n459), .A2(n1300), .B1(n462), .B2(n4020), .ZN(n2401) );
  OAI211_X1 U2718 ( .C1(n527), .C2(n465), .A(n2402), .B(n2403), .ZN(n2397) );
  AOI221_X1 U2719 ( .B1(n468), .B2(n1159), .C1(n471), .C2(n4148), .A(n2404), 
        .ZN(n2403) );
  OAI22_X1 U2720 ( .A1(n623), .A2(n474), .B1(n1620), .B2(n477), .ZN(n2404) );
  AOI22_X1 U2721 ( .A1(n480), .A2(n4180), .B1(n483), .B2(n1057), .ZN(n2402) );
  NAND4_X1 U2722 ( .A1(n2405), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n2396)
         );
  AOI221_X1 U2723 ( .B1(n486), .B2(n4212), .C1(n489), .C2(n4244), .A(n2409), 
        .ZN(n2408) );
  OAI22_X1 U2724 ( .A1(n399), .A2(n492), .B1(n367), .B2(n495), .ZN(n2409) );
  AOI221_X1 U2725 ( .B1(n498), .B2(n4276), .C1(n501), .C2(n4308), .A(n2410), 
        .ZN(n2407) );
  OAI22_X1 U2726 ( .A1(n271), .A2(n504), .B1(n239), .B2(n25), .ZN(n2410) );
  AOI221_X1 U2727 ( .B1(n507), .B2(n780), .C1(n510), .C2(n814), .A(n2411), 
        .ZN(n2406) );
  OAI22_X1 U2728 ( .A1(n1628), .A2(n513), .B1(n1629), .B2(n516), .ZN(n2411) );
  AOI221_X1 U2729 ( .B1(n551), .B2(n741), .C1(n554), .C2(n3956), .A(n2412), 
        .ZN(n2405) );
  OAI22_X1 U2730 ( .A1(n1631), .A2(n557), .B1(n1632), .B2(n560), .ZN(n2412) );
  OAI222_X1 U2731 ( .A1(n582), .A2(n432), .B1(n2413), .B2(n435), .C1(n3891), 
        .C2(n438), .ZN(n2526) );
  NOR4_X1 U2732 ( .A1(n2414), .A2(n2415), .A3(n2416), .A4(n2417), .ZN(n2413)
         );
  OAI221_X1 U2733 ( .B1(n848), .B2(n441), .C1(n1638), .C2(n444), .A(n2418), 
        .ZN(n2417) );
  AOI22_X1 U2734 ( .A1(n447), .A2(n4051), .B1(n450), .B2(n1199), .ZN(n2418) );
  OAI221_X1 U2735 ( .B1(n1640), .B2(n453), .C1(n944), .C2(n456), .A(n2419), 
        .ZN(n2416) );
  AOI22_X1 U2736 ( .A1(n459), .A2(n1301), .B1(n462), .B2(n4019), .ZN(n2419) );
  OAI211_X1 U2737 ( .C1(n528), .C2(n465), .A(n2420), .B(n2421), .ZN(n2415) );
  AOI221_X1 U2738 ( .B1(n468), .B2(n1160), .C1(n471), .C2(n4147), .A(n2422), 
        .ZN(n2421) );
  OAI22_X1 U2739 ( .A1(n624), .A2(n475), .B1(n1645), .B2(n477), .ZN(n2422) );
  AOI22_X1 U2740 ( .A1(n480), .A2(n4179), .B1(n483), .B2(n1058), .ZN(n2420) );
  NAND4_X1 U2741 ( .A1(n2423), .A2(n2426), .A3(n2425), .A4(n2424), .ZN(n2414)
         );
  AOI221_X1 U2742 ( .B1(n486), .B2(n4211), .C1(n489), .C2(n4243), .A(n2427), 
        .ZN(n2426) );
  OAI22_X1 U2743 ( .A1(n400), .A2(n492), .B1(n368), .B2(n495), .ZN(n2427) );
  AOI221_X1 U2744 ( .B1(n498), .B2(n4275), .C1(n501), .C2(n4307), .A(n2428), 
        .ZN(n2425) );
  OAI22_X1 U2745 ( .A1(n272), .A2(n504), .B1(n240), .B2(n24), .ZN(n2428) );
  AOI221_X1 U2746 ( .B1(n507), .B2(n781), .C1(n510), .C2(n815), .A(n2429), 
        .ZN(n2424) );
  OAI22_X1 U2747 ( .A1(n1653), .A2(n513), .B1(n1654), .B2(n516), .ZN(n2429) );
  AOI221_X1 U2748 ( .B1(n551), .B2(n742), .C1(n554), .C2(n3955), .A(n2430), 
        .ZN(n2423) );
  OAI22_X1 U2749 ( .A1(n1656), .A2(n557), .B1(n1657), .B2(n560), .ZN(n2430) );
  OAI222_X1 U2750 ( .A1(n581), .A2(n432), .B1(n2431), .B2(n435), .C1(n3890), 
        .C2(n438), .ZN(n2525) );
  NOR4_X1 U2751 ( .A1(n2432), .A2(n2433), .A3(n2434), .A4(n2435), .ZN(n2431)
         );
  OAI221_X1 U2752 ( .B1(n849), .B2(n441), .C1(n1663), .C2(n444), .A(n2436), 
        .ZN(n2435) );
  AOI22_X1 U2753 ( .A1(n447), .A2(n4050), .B1(n450), .B2(n1200), .ZN(n2436) );
  OAI221_X1 U2754 ( .B1(n1665), .B2(n453), .C1(n945), .C2(n456), .A(n2437), 
        .ZN(n2434) );
  AOI22_X1 U2755 ( .A1(n459), .A2(n1302), .B1(n462), .B2(n4018), .ZN(n2437) );
  OAI211_X1 U2756 ( .C1(n529), .C2(n465), .A(n2438), .B(n2439), .ZN(n2433) );
  AOI221_X1 U2757 ( .B1(n468), .B2(n1161), .C1(n471), .C2(n4146), .A(n2440), 
        .ZN(n2439) );
  OAI22_X1 U2758 ( .A1(n625), .A2(n473), .B1(n1670), .B2(n477), .ZN(n2440) );
  AOI22_X1 U2759 ( .A1(n480), .A2(n4178), .B1(n483), .B2(n1059), .ZN(n2438) );
  NAND4_X1 U2760 ( .A1(n2441), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n2432)
         );
  AOI221_X1 U2761 ( .B1(n486), .B2(n4210), .C1(n489), .C2(n4242), .A(n2445), 
        .ZN(n2444) );
  OAI22_X1 U2762 ( .A1(n401), .A2(n492), .B1(n369), .B2(n495), .ZN(n2445) );
  AOI221_X1 U2763 ( .B1(n498), .B2(n4274), .C1(n501), .C2(n4306), .A(n2446), 
        .ZN(n2443) );
  OAI22_X1 U2764 ( .A1(n273), .A2(n504), .B1(n241), .B2(n25), .ZN(n2446) );
  AOI221_X1 U2765 ( .B1(n507), .B2(n782), .C1(n510), .C2(n816), .A(n2447), 
        .ZN(n2442) );
  OAI22_X1 U2766 ( .A1(n1678), .A2(n513), .B1(n1679), .B2(n516), .ZN(n2447) );
  AOI221_X1 U2767 ( .B1(n551), .B2(n743), .C1(n554), .C2(n3954), .A(n2448), 
        .ZN(n2441) );
  OAI22_X1 U2768 ( .A1(n1681), .A2(n557), .B1(n1682), .B2(n560), .ZN(n2448) );
  OAI222_X1 U2769 ( .A1(n580), .A2(n432), .B1(n2449), .B2(n435), .C1(n3889), 
        .C2(n438), .ZN(n2524) );
  NOR4_X1 U2770 ( .A1(n2450), .A2(n2451), .A3(n2452), .A4(n2453), .ZN(n2449)
         );
  OAI221_X1 U2771 ( .B1(n850), .B2(n441), .C1(n1688), .C2(n444), .A(n2454), 
        .ZN(n2453) );
  AOI22_X1 U2772 ( .A1(n447), .A2(n4049), .B1(n450), .B2(n1201), .ZN(n2454) );
  OAI221_X1 U2773 ( .B1(n1690), .B2(n453), .C1(n946), .C2(n456), .A(n2455), 
        .ZN(n2452) );
  AOI22_X1 U2774 ( .A1(n459), .A2(n1303), .B1(n462), .B2(n4017), .ZN(n2455) );
  OAI211_X1 U2775 ( .C1(n530), .C2(n465), .A(n2456), .B(n2457), .ZN(n2451) );
  AOI221_X1 U2776 ( .B1(n468), .B2(n1162), .C1(n471), .C2(n4145), .A(n2458), 
        .ZN(n2457) );
  OAI22_X1 U2777 ( .A1(n626), .A2(n28), .B1(n1695), .B2(n477), .ZN(n2458) );
  AOI22_X1 U2778 ( .A1(n480), .A2(n4177), .B1(n483), .B2(n1060), .ZN(n2456) );
  NAND4_X1 U2779 ( .A1(n2459), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n2450)
         );
  AOI221_X1 U2780 ( .B1(n486), .B2(n4209), .C1(n489), .C2(n4241), .A(n2463), 
        .ZN(n2462) );
  OAI22_X1 U2781 ( .A1(n402), .A2(n492), .B1(n370), .B2(n495), .ZN(n2463) );
  AOI221_X1 U2782 ( .B1(n498), .B2(n4273), .C1(n501), .C2(n4305), .A(n2464), 
        .ZN(n2461) );
  OAI22_X1 U2783 ( .A1(n274), .A2(n504), .B1(n242), .B2(n24), .ZN(n2464) );
  AOI221_X1 U2784 ( .B1(n507), .B2(n783), .C1(n510), .C2(n817), .A(n2465), 
        .ZN(n2460) );
  OAI22_X1 U2785 ( .A1(n1703), .A2(n513), .B1(n1704), .B2(n516), .ZN(n2465) );
  AOI221_X1 U2786 ( .B1(n551), .B2(n744), .C1(n554), .C2(n3953), .A(n2466), 
        .ZN(n2459) );
  OAI22_X1 U2787 ( .A1(n1706), .A2(n557), .B1(n1707), .B2(n560), .ZN(n2466) );
  OAI222_X1 U2788 ( .A1(n579), .A2(n432), .B1(n2467), .B2(n435), .C1(n3888), 
        .C2(n438), .ZN(n2523) );
  OAI221_X1 U2789 ( .B1(n851), .B2(n441), .C1(n1713), .C2(n444), .A(n2472), 
        .ZN(n2471) );
  AOI22_X1 U2790 ( .A1(n447), .A2(n4048), .B1(n450), .B2(n1202), .ZN(n2472) );
  OAI221_X1 U2791 ( .B1(n1715), .B2(n453), .C1(n947), .C2(n456), .A(n2473), 
        .ZN(n2470) );
  AOI22_X1 U2792 ( .A1(n459), .A2(n1304), .B1(n462), .B2(n4016), .ZN(n2473) );
  OAI211_X1 U2793 ( .C1(n531), .C2(n465), .A(n2474), .B(n2475), .ZN(n2469) );
  AOI221_X1 U2794 ( .B1(n468), .B2(n1163), .C1(n471), .C2(n4144), .A(n2476), 
        .ZN(n2475) );
  OAI22_X1 U2795 ( .A1(n627), .A2(n27), .B1(n1720), .B2(n476), .ZN(n2476) );
  AOI22_X1 U2796 ( .A1(n480), .A2(n4176), .B1(n483), .B2(n1061), .ZN(n2474) );
  NAND4_X1 U2797 ( .A1(n2477), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n2468)
         );
  AOI221_X1 U2798 ( .B1(n486), .B2(n4208), .C1(n489), .C2(n4240), .A(n2481), 
        .ZN(n2480) );
  OAI22_X1 U2799 ( .A1(n403), .A2(n492), .B1(n371), .B2(n495), .ZN(n2481) );
  AOI221_X1 U2800 ( .B1(n498), .B2(n4272), .C1(n501), .C2(n4304), .A(n2482), 
        .ZN(n2479) );
  OAI22_X1 U2801 ( .A1(n275), .A2(n504), .B1(n243), .B2(n24), .ZN(n2482) );
  AOI221_X1 U2802 ( .B1(n507), .B2(n784), .C1(n510), .C2(n818), .A(n2483), 
        .ZN(n2478) );
  OAI22_X1 U2803 ( .A1(n1728), .A2(n513), .B1(n1729), .B2(n516), .ZN(n2483) );
  AOI221_X1 U2804 ( .B1(n551), .B2(n745), .C1(n554), .C2(n3952), .A(n2484), 
        .ZN(n2477) );
  OAI22_X1 U2805 ( .A1(n1731), .A2(n557), .B1(n1732), .B2(n560), .ZN(n2484) );
  OAI222_X1 U2806 ( .A1(n578), .A2(n432), .B1(n2485), .B2(n435), .C1(n3887), 
        .C2(n438), .ZN(n2522) );
  OAI221_X1 U2807 ( .B1(n852), .B2(n441), .C1(n1738), .C2(n444), .A(n2490), 
        .ZN(n2489) );
  AOI22_X1 U2808 ( .A1(n447), .A2(n4047), .B1(n450), .B2(n1203), .ZN(n2490) );
  OAI221_X1 U2809 ( .B1(n1740), .B2(n453), .C1(n948), .C2(n456), .A(n2491), 
        .ZN(n2488) );
  AOI22_X1 U2810 ( .A1(n459), .A2(n1305), .B1(n462), .B2(n4015), .ZN(n2491) );
  OAI211_X1 U2811 ( .C1(n532), .C2(n465), .A(n2492), .B(n2493), .ZN(n2487) );
  AOI221_X1 U2812 ( .B1(n468), .B2(n1164), .C1(n471), .C2(n4143), .A(n2494), 
        .ZN(n2493) );
  OAI22_X1 U2813 ( .A1(n628), .A2(n27), .B1(n1745), .B2(n478), .ZN(n2494) );
  AOI22_X1 U2814 ( .A1(n480), .A2(n4175), .B1(n483), .B2(n1062), .ZN(n2492) );
  NAND4_X1 U2815 ( .A1(n2495), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n2486)
         );
  AOI221_X1 U2816 ( .B1(n486), .B2(n4207), .C1(n489), .C2(n4239), .A(n2499), 
        .ZN(n2498) );
  OAI22_X1 U2817 ( .A1(n404), .A2(n492), .B1(n372), .B2(n495), .ZN(n2499) );
  AOI221_X1 U2818 ( .B1(n498), .B2(n4271), .C1(n501), .C2(n4303), .A(n2500), 
        .ZN(n2497) );
  OAI22_X1 U2819 ( .A1(n276), .A2(n504), .B1(n244), .B2(n25), .ZN(n2500) );
  AOI221_X1 U2820 ( .B1(n507), .B2(n785), .C1(n510), .C2(n819), .A(n2501), 
        .ZN(n2496) );
  OAI22_X1 U2821 ( .A1(n1753), .A2(n513), .B1(n1754), .B2(n516), .ZN(n2501) );
  AOI221_X1 U2822 ( .B1(n551), .B2(n746), .C1(n554), .C2(n3951), .A(n2502), 
        .ZN(n2495) );
  OAI22_X1 U2823 ( .A1(n1756), .A2(n557), .B1(n1757), .B2(n560), .ZN(n2502) );
  OAI222_X1 U2824 ( .A1(n577), .A2(n432), .B1(n2503), .B2(n435), .C1(n3886), 
        .C2(n438), .ZN(n2521) );
  OAI221_X1 U2825 ( .B1(n853), .B2(n441), .C1(n1763), .C2(n444), .A(n3564), 
        .ZN(n3563) );
  AOI22_X1 U2826 ( .A1(n447), .A2(n4046), .B1(n450), .B2(n1204), .ZN(n3564) );
  OAI221_X1 U2827 ( .B1(n1765), .B2(n453), .C1(n949), .C2(n456), .A(n3565), 
        .ZN(n3562) );
  AOI22_X1 U2828 ( .A1(n459), .A2(n1306), .B1(n462), .B2(n4014), .ZN(n3565) );
  OAI211_X1 U2829 ( .C1(n533), .C2(n465), .A(n3566), .B(n3567), .ZN(n2505) );
  AOI221_X1 U2830 ( .B1(n468), .B2(n1165), .C1(n471), .C2(n4142), .A(n3568), 
        .ZN(n3567) );
  OAI22_X1 U2831 ( .A1(n629), .A2(n475), .B1(n1770), .B2(n476), .ZN(n3568) );
  AOI22_X1 U2832 ( .A1(n480), .A2(n4174), .B1(n483), .B2(n1063), .ZN(n3566) );
  NAND4_X1 U2833 ( .A1(n3569), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n2504)
         );
  AOI221_X1 U2834 ( .B1(n486), .B2(n4206), .C1(n489), .C2(n4238), .A(n3573), 
        .ZN(n3572) );
  OAI22_X1 U2835 ( .A1(n405), .A2(n492), .B1(n373), .B2(n495), .ZN(n3573) );
  AOI221_X1 U2836 ( .B1(n498), .B2(n4270), .C1(n501), .C2(n4302), .A(n3574), 
        .ZN(n3571) );
  OAI22_X1 U2837 ( .A1(n277), .A2(n504), .B1(n245), .B2(n24), .ZN(n3574) );
  AOI221_X1 U2838 ( .B1(n507), .B2(n786), .C1(n510), .C2(n820), .A(n3575), 
        .ZN(n3570) );
  OAI22_X1 U2839 ( .A1(n1778), .A2(n513), .B1(n1779), .B2(n516), .ZN(n3575) );
  AOI221_X1 U2840 ( .B1(n551), .B2(n747), .C1(n554), .C2(n3950), .A(n3576), 
        .ZN(n3569) );
  OAI22_X1 U2841 ( .A1(n1781), .A2(n557), .B1(n1782), .B2(n560), .ZN(n3576) );
  OAI222_X1 U2842 ( .A1(n576), .A2(n432), .B1(n3577), .B2(n435), .C1(n3885), 
        .C2(n438), .ZN(n2520) );
  OAI221_X1 U2843 ( .B1(n854), .B2(n441), .C1(n1788), .C2(n444), .A(n3582), 
        .ZN(n3581) );
  AOI22_X1 U2844 ( .A1(n447), .A2(n4045), .B1(n450), .B2(n1205), .ZN(n3582) );
  OAI221_X1 U2845 ( .B1(n1790), .B2(n453), .C1(n950), .C2(n456), .A(n3583), 
        .ZN(n3580) );
  AOI22_X1 U2846 ( .A1(n459), .A2(n1307), .B1(n462), .B2(n4013), .ZN(n3583) );
  OAI211_X1 U2847 ( .C1(n534), .C2(n465), .A(n3584), .B(n3585), .ZN(n3579) );
  AOI221_X1 U2848 ( .B1(n468), .B2(n1166), .C1(n471), .C2(n4141), .A(n3586), 
        .ZN(n3585) );
  OAI22_X1 U2849 ( .A1(n630), .A2(n473), .B1(n1795), .B2(n478), .ZN(n3586) );
  AOI22_X1 U2850 ( .A1(n480), .A2(n4173), .B1(n483), .B2(n1064), .ZN(n3584) );
  NAND4_X1 U2851 ( .A1(n3587), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3578)
         );
  AOI221_X1 U2852 ( .B1(n486), .B2(n4205), .C1(n489), .C2(n4237), .A(n3591), 
        .ZN(n3590) );
  OAI22_X1 U2853 ( .A1(n406), .A2(n492), .B1(n374), .B2(n495), .ZN(n3591) );
  AOI221_X1 U2854 ( .B1(n498), .B2(n4269), .C1(n501), .C2(n4301), .A(n3592), 
        .ZN(n3589) );
  OAI22_X1 U2855 ( .A1(n278), .A2(n504), .B1(n246), .B2(n25), .ZN(n3592) );
  AOI221_X1 U2856 ( .B1(n507), .B2(n787), .C1(n510), .C2(n821), .A(n3593), 
        .ZN(n3588) );
  OAI22_X1 U2857 ( .A1(n1803), .A2(n513), .B1(n1804), .B2(n516), .ZN(n3593) );
  AOI221_X1 U2858 ( .B1(n551), .B2(n748), .C1(n554), .C2(n3949), .A(n3594), 
        .ZN(n3587) );
  OAI22_X1 U2859 ( .A1(n1806), .A2(n557), .B1(n1807), .B2(n560), .ZN(n3594) );
  OAI222_X1 U2860 ( .A1(n575), .A2(n432), .B1(n3595), .B2(n435), .C1(n3884), 
        .C2(n438), .ZN(n2519) );
  OAI221_X1 U2861 ( .B1(n855), .B2(n441), .C1(n1813), .C2(n444), .A(n3600), 
        .ZN(n3599) );
  AOI22_X1 U2862 ( .A1(n447), .A2(n4044), .B1(n450), .B2(n1206), .ZN(n3600) );
  OAI221_X1 U2863 ( .B1(n1815), .B2(n453), .C1(n951), .C2(n456), .A(n3601), 
        .ZN(n3598) );
  AOI22_X1 U2864 ( .A1(n459), .A2(n1308), .B1(n462), .B2(n4012), .ZN(n3601) );
  OAI211_X1 U2865 ( .C1(n535), .C2(n465), .A(n3602), .B(n3603), .ZN(n3597) );
  AOI221_X1 U2866 ( .B1(n468), .B2(n1167), .C1(n471), .C2(n4140), .A(n3604), 
        .ZN(n3603) );
  OAI22_X1 U2867 ( .A1(n631), .A2(n475), .B1(n1820), .B2(n476), .ZN(n3604) );
  AOI22_X1 U2868 ( .A1(n480), .A2(n4172), .B1(n483), .B2(n1065), .ZN(n3602) );
  NAND4_X1 U2869 ( .A1(n3605), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3596)
         );
  AOI221_X1 U2870 ( .B1(n486), .B2(n4204), .C1(n489), .C2(n4236), .A(n3609), 
        .ZN(n3608) );
  OAI22_X1 U2871 ( .A1(n407), .A2(n492), .B1(n375), .B2(n495), .ZN(n3609) );
  AOI221_X1 U2872 ( .B1(n498), .B2(n4268), .C1(n501), .C2(n4300), .A(n3610), 
        .ZN(n3607) );
  OAI22_X1 U2873 ( .A1(n279), .A2(n504), .B1(n247), .B2(n24), .ZN(n3610) );
  AOI221_X1 U2874 ( .B1(n507), .B2(n788), .C1(n510), .C2(n822), .A(n3611), 
        .ZN(n3606) );
  OAI22_X1 U2875 ( .A1(n1828), .A2(n513), .B1(n1829), .B2(n516), .ZN(n3611) );
  AOI221_X1 U2876 ( .B1(n551), .B2(n749), .C1(n554), .C2(n3948), .A(n3612), 
        .ZN(n3605) );
  OAI22_X1 U2877 ( .A1(n1831), .A2(n557), .B1(n1832), .B2(n560), .ZN(n3612) );
  OAI222_X1 U2878 ( .A1(n574), .A2(n432), .B1(n3613), .B2(n435), .C1(n3883), 
        .C2(n438), .ZN(n2518) );
  OAI221_X1 U2879 ( .B1(n856), .B2(n441), .C1(n1838), .C2(n444), .A(n3618), 
        .ZN(n3617) );
  AOI22_X1 U2880 ( .A1(n447), .A2(n4043), .B1(n450), .B2(n1207), .ZN(n3618) );
  OAI221_X1 U2881 ( .B1(n1840), .B2(n453), .C1(n952), .C2(n456), .A(n3619), 
        .ZN(n3616) );
  AOI22_X1 U2882 ( .A1(n459), .A2(n1309), .B1(n462), .B2(n4011), .ZN(n3619) );
  OAI211_X1 U2883 ( .C1(n536), .C2(n465), .A(n3620), .B(n3621), .ZN(n3615) );
  AOI221_X1 U2884 ( .B1(n468), .B2(n1168), .C1(n471), .C2(n4139), .A(n3622), 
        .ZN(n3621) );
  OAI22_X1 U2885 ( .A1(n632), .A2(n473), .B1(n1845), .B2(n478), .ZN(n3622) );
  AOI22_X1 U2886 ( .A1(n480), .A2(n4171), .B1(n483), .B2(n1066), .ZN(n3620) );
  NAND4_X1 U2887 ( .A1(n3623), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3614)
         );
  AOI221_X1 U2888 ( .B1(n486), .B2(n4203), .C1(n489), .C2(n4235), .A(n3627), 
        .ZN(n3626) );
  OAI22_X1 U2889 ( .A1(n408), .A2(n492), .B1(n376), .B2(n495), .ZN(n3627) );
  AOI221_X1 U2890 ( .B1(n498), .B2(n4267), .C1(n501), .C2(n4299), .A(n3628), 
        .ZN(n3625) );
  OAI22_X1 U2891 ( .A1(n280), .A2(n504), .B1(n248), .B2(n25), .ZN(n3628) );
  AOI221_X1 U2892 ( .B1(n507), .B2(n789), .C1(n510), .C2(n823), .A(n3629), 
        .ZN(n3624) );
  OAI22_X1 U2893 ( .A1(n1853), .A2(n513), .B1(n1854), .B2(n516), .ZN(n3629) );
  AOI221_X1 U2894 ( .B1(n551), .B2(n750), .C1(n554), .C2(n3947), .A(n3630), 
        .ZN(n3623) );
  OAI22_X1 U2895 ( .A1(n1856), .A2(n557), .B1(n1857), .B2(n560), .ZN(n3630) );
  OAI222_X1 U2896 ( .A1(n573), .A2(n431), .B1(n3631), .B2(n434), .C1(n3882), 
        .C2(n438), .ZN(n2517) );
  NOR4_X1 U2897 ( .A1(n3632), .A2(n3633), .A3(n3634), .A4(n3635), .ZN(n3631)
         );
  OAI221_X1 U2898 ( .B1(n857), .B2(n440), .C1(n1863), .C2(n443), .A(n3636), 
        .ZN(n3635) );
  AOI22_X1 U2899 ( .A1(n446), .A2(n4042), .B1(n449), .B2(n1208), .ZN(n3636) );
  OAI221_X1 U2900 ( .B1(n1865), .B2(n452), .C1(n953), .C2(n455), .A(n3637), 
        .ZN(n3634) );
  AOI22_X1 U2901 ( .A1(n458), .A2(n1310), .B1(n461), .B2(n4010), .ZN(n3637) );
  OAI211_X1 U2902 ( .C1(n537), .C2(n464), .A(n3638), .B(n3639), .ZN(n3633) );
  AOI221_X1 U2903 ( .B1(n467), .B2(n1169), .C1(n470), .C2(n4138), .A(n3640), 
        .ZN(n3639) );
  OAI22_X1 U2904 ( .A1(n633), .A2(n474), .B1(n1870), .B2(n477), .ZN(n3640) );
  AOI22_X1 U2905 ( .A1(n479), .A2(n4170), .B1(n482), .B2(n1067), .ZN(n3638) );
  NAND4_X1 U2906 ( .A1(n3641), .A2(n3642), .A3(n3643), .A4(n3644), .ZN(n3632)
         );
  AOI221_X1 U2907 ( .B1(n485), .B2(n4202), .C1(n488), .C2(n4234), .A(n3645), 
        .ZN(n3644) );
  OAI22_X1 U2908 ( .A1(n409), .A2(n491), .B1(n377), .B2(n494), .ZN(n3645) );
  AOI221_X1 U2909 ( .B1(n497), .B2(n4266), .C1(n500), .C2(n4298), .A(n3646), 
        .ZN(n3643) );
  OAI22_X1 U2910 ( .A1(n281), .A2(n503), .B1(n249), .B2(n24), .ZN(n3646) );
  OAI22_X1 U2911 ( .A1(n1878), .A2(n512), .B1(n1879), .B2(n515), .ZN(n3647) );
  AOI221_X1 U2912 ( .B1(n550), .B2(n751), .C1(n553), .C2(n3946), .A(n3648), 
        .ZN(n3641) );
  OAI22_X1 U2913 ( .A1(n1881), .A2(n556), .B1(n1882), .B2(n559), .ZN(n3648) );
  OAI222_X1 U2914 ( .A1(n572), .A2(n431), .B1(n3649), .B2(n434), .C1(n3881), 
        .C2(n438), .ZN(n2516) );
  NOR4_X1 U2915 ( .A1(n3650), .A2(n3651), .A3(n3652), .A4(n3653), .ZN(n3649)
         );
  OAI221_X1 U2916 ( .B1(n858), .B2(n440), .C1(n1888), .C2(n443), .A(n3654), 
        .ZN(n3653) );
  AOI22_X1 U2917 ( .A1(n446), .A2(n4041), .B1(n449), .B2(n1209), .ZN(n3654) );
  OAI221_X1 U2918 ( .B1(n1890), .B2(n452), .C1(n954), .C2(n455), .A(n3655), 
        .ZN(n3652) );
  AOI22_X1 U2919 ( .A1(n458), .A2(n1311), .B1(n461), .B2(n4009), .ZN(n3655) );
  OAI211_X1 U2920 ( .C1(n538), .C2(n464), .A(n3656), .B(n3657), .ZN(n3651) );
  AOI221_X1 U2921 ( .B1(n467), .B2(n1170), .C1(n470), .C2(n4137), .A(n3658), 
        .ZN(n3657) );
  OAI22_X1 U2922 ( .A1(n634), .A2(n474), .B1(n1895), .B2(n477), .ZN(n3658) );
  AOI22_X1 U2923 ( .A1(n479), .A2(n4169), .B1(n482), .B2(n1068), .ZN(n3656) );
  NAND4_X1 U2924 ( .A1(n3659), .A2(n3660), .A3(n3661), .A4(n3662), .ZN(n3650)
         );
  AOI221_X1 U2925 ( .B1(n485), .B2(n4201), .C1(n488), .C2(n4233), .A(n3663), 
        .ZN(n3662) );
  OAI22_X1 U2926 ( .A1(n410), .A2(n491), .B1(n378), .B2(n494), .ZN(n3663) );
  AOI221_X1 U2927 ( .B1(n497), .B2(n4265), .C1(n500), .C2(n4297), .A(n3664), 
        .ZN(n3661) );
  OAI22_X1 U2928 ( .A1(n282), .A2(n503), .B1(n250), .B2(n25), .ZN(n3664) );
  OAI22_X1 U2929 ( .A1(n1903), .A2(n512), .B1(n1904), .B2(n515), .ZN(n3665) );
  AOI221_X1 U2930 ( .B1(n550), .B2(n752), .C1(n553), .C2(n3945), .A(n3666), 
        .ZN(n3659) );
  OAI22_X1 U2931 ( .A1(n1906), .A2(n556), .B1(n1907), .B2(n559), .ZN(n3666) );
  OAI222_X1 U2932 ( .A1(n571), .A2(n431), .B1(n3667), .B2(n434), .C1(n3880), 
        .C2(n437), .ZN(n2515) );
  OAI221_X1 U2933 ( .B1(n859), .B2(n440), .C1(n1913), .C2(n443), .A(n3672), 
        .ZN(n3671) );
  AOI22_X1 U2934 ( .A1(n446), .A2(n4040), .B1(n449), .B2(n1210), .ZN(n3672) );
  OAI221_X1 U2935 ( .B1(n1915), .B2(n452), .C1(n955), .C2(n455), .A(n3673), 
        .ZN(n3670) );
  AOI22_X1 U2936 ( .A1(n458), .A2(n1312), .B1(n461), .B2(n4008), .ZN(n3673) );
  OAI211_X1 U2937 ( .C1(n539), .C2(n464), .A(n3674), .B(n3675), .ZN(n3669) );
  AOI221_X1 U2938 ( .B1(n467), .B2(n1171), .C1(n470), .C2(n4136), .A(n3676), 
        .ZN(n3675) );
  OAI22_X1 U2939 ( .A1(n635), .A2(n475), .B1(n1920), .B2(n476), .ZN(n3676) );
  AOI22_X1 U2940 ( .A1(n479), .A2(n4168), .B1(n482), .B2(n1069), .ZN(n3674) );
  NAND4_X1 U2941 ( .A1(n3677), .A2(n3678), .A3(n3679), .A4(n3680), .ZN(n3668)
         );
  AOI221_X1 U2942 ( .B1(n485), .B2(n4200), .C1(n488), .C2(n4232), .A(n3681), 
        .ZN(n3680) );
  OAI22_X1 U2943 ( .A1(n411), .A2(n491), .B1(n379), .B2(n494), .ZN(n3681) );
  AOI221_X1 U2944 ( .B1(n497), .B2(n4264), .C1(n500), .C2(n4296), .A(n3682), 
        .ZN(n3679) );
  OAI22_X1 U2945 ( .A1(n283), .A2(n503), .B1(n251), .B2(n24), .ZN(n3682) );
  AOI221_X1 U2946 ( .B1(n506), .B2(n792), .C1(n509), .C2(n826), .A(n3683), 
        .ZN(n3678) );
  OAI22_X1 U2947 ( .A1(n1928), .A2(n512), .B1(n1929), .B2(n515), .ZN(n3683) );
  AOI221_X1 U2948 ( .B1(n550), .B2(n753), .C1(n553), .C2(n3944), .A(n3684), 
        .ZN(n3677) );
  OAI22_X1 U2949 ( .A1(n1931), .A2(n556), .B1(n1932), .B2(n559), .ZN(n3684) );
  OAI222_X1 U2950 ( .A1(n570), .A2(n431), .B1(n3685), .B2(n434), .C1(n3879), 
        .C2(n437), .ZN(n2514) );
  OAI221_X1 U2951 ( .B1(n860), .B2(n440), .C1(n1938), .C2(n443), .A(n3690), 
        .ZN(n3689) );
  AOI22_X1 U2952 ( .A1(n446), .A2(n4039), .B1(n449), .B2(n1211), .ZN(n3690) );
  OAI221_X1 U2953 ( .B1(n1940), .B2(n452), .C1(n956), .C2(n455), .A(n3691), 
        .ZN(n3688) );
  AOI22_X1 U2954 ( .A1(n458), .A2(n1313), .B1(n461), .B2(n4007), .ZN(n3691) );
  OAI211_X1 U2955 ( .C1(n540), .C2(n464), .A(n3692), .B(n3693), .ZN(n3687) );
  AOI221_X1 U2956 ( .B1(n467), .B2(n1172), .C1(n470), .C2(n4135), .A(n3694), 
        .ZN(n3693) );
  OAI22_X1 U2957 ( .A1(n636), .A2(n475), .B1(n1945), .B2(n478), .ZN(n3694) );
  AOI22_X1 U2958 ( .A1(n479), .A2(n4167), .B1(n482), .B2(n1070), .ZN(n3692) );
  NAND4_X1 U2959 ( .A1(n3695), .A2(n3696), .A3(n3697), .A4(n3698), .ZN(n3686)
         );
  AOI221_X1 U2960 ( .B1(n485), .B2(n4199), .C1(n488), .C2(n4231), .A(n3699), 
        .ZN(n3698) );
  OAI22_X1 U2961 ( .A1(n412), .A2(n491), .B1(n380), .B2(n494), .ZN(n3699) );
  AOI221_X1 U2962 ( .B1(n497), .B2(n4263), .C1(n500), .C2(n4295), .A(n3700), 
        .ZN(n3697) );
  OAI22_X1 U2963 ( .A1(n284), .A2(n503), .B1(n252), .B2(n25), .ZN(n3700) );
  OAI22_X1 U2964 ( .A1(n1953), .A2(n512), .B1(n1954), .B2(n515), .ZN(n3701) );
  AOI221_X1 U2965 ( .B1(n550), .B2(n754), .C1(n553), .C2(n3943), .A(n3702), 
        .ZN(n3695) );
  OAI22_X1 U2966 ( .A1(n1956), .A2(n556), .B1(n1957), .B2(n559), .ZN(n3702) );
  OAI222_X1 U2967 ( .A1(n569), .A2(n431), .B1(n3703), .B2(n434), .C1(n3878), 
        .C2(n437), .ZN(n2513) );
  NOR4_X1 U2968 ( .A1(n3704), .A2(n3705), .A3(n3706), .A4(n3707), .ZN(n3703)
         );
  OAI221_X1 U2969 ( .B1(n861), .B2(n440), .C1(n1963), .C2(n443), .A(n3708), 
        .ZN(n3707) );
  AOI22_X1 U2970 ( .A1(n446), .A2(n4038), .B1(n449), .B2(n1212), .ZN(n3708) );
  OAI221_X1 U2971 ( .B1(n1965), .B2(n452), .C1(n957), .C2(n455), .A(n3709), 
        .ZN(n3706) );
  AOI22_X1 U2972 ( .A1(n458), .A2(n1314), .B1(n461), .B2(n4006), .ZN(n3709) );
  OAI211_X1 U2973 ( .C1(n541), .C2(n464), .A(n3710), .B(n3711), .ZN(n3705) );
  AOI221_X1 U2974 ( .B1(n467), .B2(n1173), .C1(n470), .C2(n4134), .A(n3712), 
        .ZN(n3711) );
  OAI22_X1 U2975 ( .A1(n637), .A2(n474), .B1(n1970), .B2(n477), .ZN(n3712) );
  AOI22_X1 U2976 ( .A1(n479), .A2(n4166), .B1(n482), .B2(n1071), .ZN(n3710) );
  NAND4_X1 U2977 ( .A1(n3713), .A2(n3714), .A3(n3715), .A4(n3716), .ZN(n3704)
         );
  AOI221_X1 U2978 ( .B1(n485), .B2(n4198), .C1(n488), .C2(n4230), .A(n3717), 
        .ZN(n3716) );
  OAI22_X1 U2979 ( .A1(n413), .A2(n491), .B1(n381), .B2(n494), .ZN(n3717) );
  AOI221_X1 U2980 ( .B1(n497), .B2(n4262), .C1(n500), .C2(n4294), .A(n3718), 
        .ZN(n3715) );
  OAI22_X1 U2981 ( .A1(n285), .A2(n503), .B1(n253), .B2(n24), .ZN(n3718) );
  OAI22_X1 U2982 ( .A1(n1978), .A2(n512), .B1(n1979), .B2(n515), .ZN(n3719) );
  AOI221_X1 U2983 ( .B1(n550), .B2(n755), .C1(n553), .C2(n3942), .A(n3720), 
        .ZN(n3713) );
  OAI22_X1 U2984 ( .A1(n1981), .A2(n556), .B1(n1982), .B2(n559), .ZN(n3720) );
  OAI222_X1 U2985 ( .A1(n568), .A2(n431), .B1(n3721), .B2(n434), .C1(n3877), 
        .C2(n437), .ZN(n2512) );
  OAI221_X1 U2986 ( .B1(n862), .B2(n440), .C1(n1988), .C2(n443), .A(n3726), 
        .ZN(n3725) );
  AOI22_X1 U2987 ( .A1(n446), .A2(n4037), .B1(n449), .B2(n1213), .ZN(n3726) );
  OAI221_X1 U2988 ( .B1(n1990), .B2(n452), .C1(n958), .C2(n455), .A(n3727), 
        .ZN(n3724) );
  AOI22_X1 U2989 ( .A1(n458), .A2(n1315), .B1(n461), .B2(n4005), .ZN(n3727) );
  OAI211_X1 U2990 ( .C1(n542), .C2(n464), .A(n3728), .B(n3729), .ZN(n3723) );
  AOI221_X1 U2991 ( .B1(n467), .B2(n1174), .C1(n470), .C2(n4133), .A(n3730), 
        .ZN(n3729) );
  OAI22_X1 U2992 ( .A1(n638), .A2(n28), .B1(n1995), .B2(n476), .ZN(n3730) );
  AOI22_X1 U2993 ( .A1(n479), .A2(n4165), .B1(n482), .B2(n1072), .ZN(n3728) );
  NAND4_X1 U2994 ( .A1(n3731), .A2(n3732), .A3(n3733), .A4(n3734), .ZN(n3722)
         );
  AOI221_X1 U2995 ( .B1(n485), .B2(n4197), .C1(n488), .C2(n4229), .A(n3735), 
        .ZN(n3734) );
  OAI22_X1 U2996 ( .A1(n414), .A2(n491), .B1(n382), .B2(n494), .ZN(n3735) );
  AOI221_X1 U2997 ( .B1(n497), .B2(n4261), .C1(n500), .C2(n4293), .A(n3736), 
        .ZN(n3733) );
  OAI22_X1 U2998 ( .A1(n286), .A2(n503), .B1(n254), .B2(n24), .ZN(n3736) );
  OAI22_X1 U2999 ( .A1(n2003), .A2(n512), .B1(n2004), .B2(n515), .ZN(n3737) );
  AOI221_X1 U3000 ( .B1(n550), .B2(n756), .C1(n553), .C2(n3941), .A(n3738), 
        .ZN(n3731) );
  OAI22_X1 U3001 ( .A1(n2006), .A2(n556), .B1(n2007), .B2(n559), .ZN(n3738) );
  OAI222_X1 U3002 ( .A1(n567), .A2(n431), .B1(n3739), .B2(n434), .C1(n3876), 
        .C2(n437), .ZN(n2511) );
  OAI221_X1 U3003 ( .B1(n863), .B2(n440), .C1(n2013), .C2(n443), .A(n3744), 
        .ZN(n3743) );
  AOI22_X1 U3004 ( .A1(n446), .A2(n4036), .B1(n449), .B2(n1214), .ZN(n3744) );
  OAI221_X1 U3005 ( .B1(n2015), .B2(n452), .C1(n959), .C2(n455), .A(n3745), 
        .ZN(n3742) );
  AOI22_X1 U3006 ( .A1(n458), .A2(n1316), .B1(n461), .B2(n4004), .ZN(n3745) );
  OAI211_X1 U3007 ( .C1(n543), .C2(n464), .A(n3746), .B(n3747), .ZN(n3741) );
  AOI221_X1 U3008 ( .B1(n467), .B2(n1175), .C1(n470), .C2(n4132), .A(n3748), 
        .ZN(n3747) );
  OAI22_X1 U3009 ( .A1(n639), .A2(n27), .B1(n2020), .B2(n478), .ZN(n3748) );
  AOI22_X1 U3010 ( .A1(n479), .A2(n4164), .B1(n482), .B2(n1073), .ZN(n3746) );
  NAND4_X1 U3011 ( .A1(n3749), .A2(n3750), .A3(n3751), .A4(n3752), .ZN(n3740)
         );
  AOI221_X1 U3012 ( .B1(n485), .B2(n4196), .C1(n488), .C2(n4228), .A(n3753), 
        .ZN(n3752) );
  OAI22_X1 U3013 ( .A1(n415), .A2(n491), .B1(n383), .B2(n494), .ZN(n3753) );
  AOI221_X1 U3014 ( .B1(n497), .B2(n4260), .C1(n500), .C2(n4292), .A(n3754), 
        .ZN(n3751) );
  OAI22_X1 U3015 ( .A1(n287), .A2(n503), .B1(n255), .B2(n25), .ZN(n3754) );
  OAI22_X1 U3016 ( .A1(n2028), .A2(n512), .B1(n2029), .B2(n515), .ZN(n3755) );
  AOI221_X1 U3017 ( .B1(n550), .B2(n757), .C1(n553), .C2(n3940), .A(n3756), 
        .ZN(n3749) );
  OAI22_X1 U3018 ( .A1(n2031), .A2(n556), .B1(n2032), .B2(n559), .ZN(n3756) );
  OAI222_X1 U3019 ( .A1(n566), .A2(n431), .B1(n3757), .B2(n434), .C1(n3875), 
        .C2(n437), .ZN(n2510) );
  OAI221_X1 U3020 ( .B1(n864), .B2(n440), .C1(n2038), .C2(n443), .A(n3762), 
        .ZN(n3761) );
  AOI22_X1 U3021 ( .A1(n446), .A2(n4035), .B1(n449), .B2(n1215), .ZN(n3762) );
  OAI221_X1 U3022 ( .B1(n2040), .B2(n452), .C1(n960), .C2(n455), .A(n3763), 
        .ZN(n3760) );
  AOI22_X1 U3023 ( .A1(n458), .A2(n1317), .B1(n461), .B2(n4003), .ZN(n3763) );
  OAI211_X1 U3024 ( .C1(n544), .C2(n464), .A(n3764), .B(n3765), .ZN(n3759) );
  AOI221_X1 U3025 ( .B1(n467), .B2(n1176), .C1(n470), .C2(n4131), .A(n3766), 
        .ZN(n3765) );
  OAI22_X1 U3026 ( .A1(n640), .A2(n473), .B1(n2045), .B2(n476), .ZN(n3766) );
  AOI22_X1 U3027 ( .A1(n479), .A2(n4163), .B1(n482), .B2(n1074), .ZN(n3764) );
  NAND4_X1 U3028 ( .A1(n3767), .A2(n3768), .A3(n3769), .A4(n3770), .ZN(n3758)
         );
  AOI221_X1 U3029 ( .B1(n485), .B2(n4195), .C1(n488), .C2(n4227), .A(n3771), 
        .ZN(n3770) );
  OAI22_X1 U3030 ( .A1(n416), .A2(n491), .B1(n384), .B2(n494), .ZN(n3771) );
  AOI221_X1 U3031 ( .B1(n497), .B2(n4259), .C1(n500), .C2(n4291), .A(n3772), 
        .ZN(n3769) );
  OAI22_X1 U3032 ( .A1(n288), .A2(n503), .B1(n256), .B2(n24), .ZN(n3772) );
  AOI221_X1 U3033 ( .B1(n506), .B2(n797), .C1(n509), .C2(n831), .A(n3773), 
        .ZN(n3768) );
  OAI22_X1 U3034 ( .A1(n2053), .A2(n512), .B1(n2054), .B2(n515), .ZN(n3773) );
  AOI221_X1 U3035 ( .B1(n550), .B2(n758), .C1(n553), .C2(n3939), .A(n3774), 
        .ZN(n3767) );
  OAI22_X1 U3036 ( .A1(n2056), .A2(n556), .B1(n2057), .B2(n559), .ZN(n3774) );
  OAI222_X1 U3037 ( .A1(n565), .A2(n431), .B1(n3775), .B2(n434), .C1(n3874), 
        .C2(n437), .ZN(n2509) );
  OAI221_X1 U3038 ( .B1(n865), .B2(n440), .C1(n2063), .C2(n443), .A(n3780), 
        .ZN(n3779) );
  AOI22_X1 U3039 ( .A1(n446), .A2(n4034), .B1(n449), .B2(n1216), .ZN(n3780) );
  OAI221_X1 U3040 ( .B1(n2065), .B2(n452), .C1(n961), .C2(n455), .A(n3781), 
        .ZN(n3778) );
  AOI22_X1 U3041 ( .A1(n458), .A2(n1318), .B1(n461), .B2(n4002), .ZN(n3781) );
  OAI211_X1 U3042 ( .C1(n545), .C2(n464), .A(n3782), .B(n3783), .ZN(n3777) );
  AOI221_X1 U3043 ( .B1(n467), .B2(n1177), .C1(n470), .C2(n4130), .A(n3784), 
        .ZN(n3783) );
  OAI22_X1 U3044 ( .A1(n641), .A2(n28), .B1(n2070), .B2(n478), .ZN(n3784) );
  AOI22_X1 U3045 ( .A1(n479), .A2(n4162), .B1(n482), .B2(n1075), .ZN(n3782) );
  NAND4_X1 U3046 ( .A1(n3785), .A2(n3786), .A3(n3787), .A4(n3788), .ZN(n3776)
         );
  AOI221_X1 U3047 ( .B1(n485), .B2(n4194), .C1(n488), .C2(n4226), .A(n3789), 
        .ZN(n3788) );
  OAI22_X1 U3048 ( .A1(n417), .A2(n491), .B1(n385), .B2(n494), .ZN(n3789) );
  AOI221_X1 U3049 ( .B1(n497), .B2(n4258), .C1(n500), .C2(n4290), .A(n3790), 
        .ZN(n3787) );
  OAI22_X1 U3050 ( .A1(n289), .A2(n503), .B1(n257), .B2(n25), .ZN(n3790) );
  AOI221_X1 U3051 ( .B1(n506), .B2(n798), .C1(n509), .C2(n832), .A(n3791), 
        .ZN(n3786) );
  OAI22_X1 U3052 ( .A1(n2078), .A2(n512), .B1(n2079), .B2(n515), .ZN(n3791) );
  AOI221_X1 U3053 ( .B1(n550), .B2(n759), .C1(n553), .C2(n3938), .A(n3792), 
        .ZN(n3785) );
  OAI22_X1 U3054 ( .A1(n2081), .A2(n556), .B1(n2082), .B2(n559), .ZN(n3792) );
  OAI222_X1 U3055 ( .A1(n564), .A2(n431), .B1(n3793), .B2(n434), .C1(n3873), 
        .C2(n437), .ZN(n2508) );
  OAI221_X1 U3056 ( .B1(n866), .B2(n440), .C1(n2088), .C2(n443), .A(n3798), 
        .ZN(n3797) );
  AOI22_X1 U3057 ( .A1(n446), .A2(n4033), .B1(n449), .B2(n1217), .ZN(n3798) );
  OAI221_X1 U3058 ( .B1(n2090), .B2(n452), .C1(n962), .C2(n455), .A(n3799), 
        .ZN(n3796) );
  AOI22_X1 U3059 ( .A1(n458), .A2(n1319), .B1(n461), .B2(n4001), .ZN(n3799) );
  OAI211_X1 U3060 ( .C1(n546), .C2(n464), .A(n3800), .B(n3801), .ZN(n3795) );
  AOI221_X1 U3061 ( .B1(n467), .B2(n1178), .C1(n470), .C2(n4129), .A(n3802), 
        .ZN(n3801) );
  OAI22_X1 U3062 ( .A1(n642), .A2(n27), .B1(n2095), .B2(n476), .ZN(n3802) );
  AOI22_X1 U3063 ( .A1(n479), .A2(n4161), .B1(n482), .B2(n1076), .ZN(n3800) );
  NAND4_X1 U3064 ( .A1(n3803), .A2(n3804), .A3(n3805), .A4(n3806), .ZN(n3794)
         );
  AOI221_X1 U3065 ( .B1(n485), .B2(n4193), .C1(n488), .C2(n4225), .A(n3807), 
        .ZN(n3806) );
  OAI22_X1 U3066 ( .A1(n418), .A2(n491), .B1(n386), .B2(n494), .ZN(n3807) );
  AOI221_X1 U3067 ( .B1(n497), .B2(n4257), .C1(n500), .C2(n4289), .A(n3808), 
        .ZN(n3805) );
  OAI22_X1 U3068 ( .A1(n290), .A2(n503), .B1(n258), .B2(n24), .ZN(n3808) );
  OAI22_X1 U3069 ( .A1(n2103), .A2(n512), .B1(n2104), .B2(n515), .ZN(n3809) );
  AOI221_X1 U3070 ( .B1(n550), .B2(n760), .C1(n553), .C2(n3937), .A(n3810), 
        .ZN(n3803) );
  OAI22_X1 U3071 ( .A1(n2106), .A2(n556), .B1(n2107), .B2(n559), .ZN(n3810) );
  OAI222_X1 U3072 ( .A1(n563), .A2(n431), .B1(n3811), .B2(n434), .C1(n3872), 
        .C2(n437), .ZN(n2507) );
  OAI221_X1 U3073 ( .B1(n867), .B2(n440), .C1(n2113), .C2(n443), .A(n3816), 
        .ZN(n3815) );
  AOI22_X1 U3074 ( .A1(n446), .A2(n4032), .B1(n449), .B2(n1218), .ZN(n3816) );
  OAI221_X1 U3075 ( .B1(n2115), .B2(n452), .C1(n963), .C2(n455), .A(n3817), 
        .ZN(n3814) );
  AOI22_X1 U3076 ( .A1(n458), .A2(n1320), .B1(n461), .B2(n4000), .ZN(n3817) );
  OAI211_X1 U3077 ( .C1(n547), .C2(n464), .A(n3818), .B(n3819), .ZN(n3813) );
  AOI221_X1 U3078 ( .B1(n467), .B2(n1179), .C1(n470), .C2(n4128), .A(n3820), 
        .ZN(n3819) );
  OAI22_X1 U3079 ( .A1(n643), .A2(n475), .B1(n2120), .B2(n478), .ZN(n3820) );
  AOI22_X1 U3080 ( .A1(n479), .A2(n4160), .B1(n482), .B2(n1077), .ZN(n3818) );
  NAND4_X1 U3081 ( .A1(n3821), .A2(n3822), .A3(n3823), .A4(n3824), .ZN(n3812)
         );
  AOI221_X1 U3082 ( .B1(n485), .B2(n4192), .C1(n488), .C2(n4224), .A(n3825), 
        .ZN(n3824) );
  OAI22_X1 U3083 ( .A1(n419), .A2(n491), .B1(n387), .B2(n494), .ZN(n3825) );
  AOI221_X1 U3084 ( .B1(n497), .B2(n4256), .C1(n500), .C2(n4288), .A(n3826), 
        .ZN(n3823) );
  OAI22_X1 U3085 ( .A1(n291), .A2(n503), .B1(n259), .B2(n25), .ZN(n3826) );
  AOI221_X1 U3086 ( .B1(n506), .B2(n800), .C1(n509), .C2(n834), .A(n3827), 
        .ZN(n3822) );
  OAI22_X1 U3087 ( .A1(n2128), .A2(n512), .B1(n2129), .B2(n515), .ZN(n3827) );
  AOI221_X1 U3088 ( .B1(n550), .B2(n761), .C1(n553), .C2(n3936), .A(n3828), 
        .ZN(n3821) );
  OAI22_X1 U3089 ( .A1(n2131), .A2(n556), .B1(n2132), .B2(n559), .ZN(n3828) );
  OAI222_X1 U3090 ( .A1(n562), .A2(n431), .B1(n3829), .B2(n434), .C1(n3871), 
        .C2(n437), .ZN(n2506) );
  NAND2_X1 U3091 ( .A1(n437), .A2(n3830), .ZN(n2183) );
  NOR4_X1 U3092 ( .A1(n3831), .A2(n3832), .A3(n3833), .A4(n3834), .ZN(n3829)
         );
  OAI221_X1 U3093 ( .B1(n868), .B2(n440), .C1(n2139), .C2(n443), .A(n3835), 
        .ZN(n3834) );
  AOI22_X1 U3094 ( .A1(n446), .A2(n4031), .B1(n449), .B2(n1219), .ZN(n3835) );
  AND2_X1 U3095 ( .A1(n3836), .A2(n3837), .ZN(n2193) );
  AND2_X1 U3096 ( .A1(n3836), .A2(n3838), .ZN(n2192) );
  NAND2_X1 U3097 ( .A1(n3839), .A2(n3840), .ZN(n2190) );
  NAND2_X1 U3098 ( .A1(n3841), .A2(n3837), .ZN(n2189) );
  OAI221_X1 U3099 ( .B1(n2147), .B2(n452), .C1(n964), .C2(n455), .A(n3842), 
        .ZN(n3833) );
  AOI22_X1 U3100 ( .A1(n458), .A2(n1321), .B1(n461), .B2(n3999), .ZN(n3842) );
  AND2_X1 U3101 ( .A1(n3841), .A2(n3838), .ZN(n2198) );
  AND2_X1 U3102 ( .A1(n3841), .A2(n3840), .ZN(n2197) );
  NAND2_X1 U3103 ( .A1(n3836), .A2(n3840), .ZN(n2195) );
  NAND2_X1 U3104 ( .A1(n3836), .A2(n113), .ZN(n2194) );
  NOR3_X1 U3105 ( .A1(n55), .A2(ADD_RS1[0]), .A3(n3844), .ZN(n3836) );
  OAI211_X1 U3106 ( .C1(n548), .C2(n464), .A(n3845), .B(n3846), .ZN(n3832) );
  OAI22_X1 U3107 ( .A1(n644), .A2(n28), .B1(n2155), .B2(n476), .ZN(n3847) );
  NAND2_X1 U3108 ( .A1(n2), .A2(n3840), .ZN(n2206) );
  NAND2_X1 U3109 ( .A1(n3848), .A2(n3843), .ZN(n2205) );
  AND2_X1 U3110 ( .A1(n3839), .A2(n3837), .ZN(n2203) );
  AND2_X1 U3111 ( .A1(n3839), .A2(n113), .ZN(n2202) );
  AOI22_X1 U3112 ( .A1(n479), .A2(n4159), .B1(n482), .B2(n1078), .ZN(n3845) );
  AND2_X1 U3113 ( .A1(n58), .A2(n3838), .ZN(n2208) );
  AND2_X1 U3114 ( .A1(n58), .A2(n3837), .ZN(n2207) );
  NOR3_X1 U3115 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[3]), .A3(n56), .ZN(n3848) );
  NAND2_X1 U3116 ( .A1(n3839), .A2(n3838), .ZN(n2199) );
  NOR3_X1 U3117 ( .A1(n83), .A2(ADD_RS1[3]), .A3(n55), .ZN(n3839) );
  NAND4_X1 U3118 ( .A1(n3849), .A2(n3850), .A3(n3851), .A4(n3852), .ZN(n3831)
         );
  AOI221_X1 U3119 ( .B1(n485), .B2(n4191), .C1(n488), .C2(n4223), .A(n3853), 
        .ZN(n3852) );
  OAI22_X1 U3120 ( .A1(n420), .A2(n491), .B1(n388), .B2(n494), .ZN(n3853) );
  NAND2_X1 U3121 ( .A1(n3843), .A2(n3854), .ZN(n2217) );
  NAND2_X1 U3122 ( .A1(n113), .A2(n3855), .ZN(n2216) );
  AND2_X1 U3123 ( .A1(n36), .A2(n3840), .ZN(n2214) );
  AND2_X1 U3124 ( .A1(n3840), .A2(n3855), .ZN(n2213) );
  AOI221_X1 U3125 ( .B1(n497), .B2(n4255), .C1(n500), .C2(n4287), .A(n3856), 
        .ZN(n3851) );
  OAI22_X1 U3126 ( .A1(n292), .A2(n503), .B1(n260), .B2(n25), .ZN(n3856) );
  NAND2_X1 U3127 ( .A1(n3838), .A2(n3854), .ZN(n2222) );
  NAND2_X1 U3128 ( .A1(n3838), .A2(n3855), .ZN(n2221) );
  AND2_X1 U3129 ( .A1(n3837), .A2(n36), .ZN(n2219) );
  NOR3_X1 U3130 ( .A1(ADD_RS1[0]), .A2(ADD_RS1[4]), .A3(n3844), .ZN(n3854) );
  AND2_X1 U3131 ( .A1(n3837), .A2(n3855), .ZN(n2218) );
  OAI22_X1 U3132 ( .A1(n2166), .A2(n512), .B1(n2167), .B2(n515), .ZN(n3857) );
  NAND2_X1 U3133 ( .A1(n3858), .A2(n3840), .ZN(n2227) );
  NAND2_X1 U3134 ( .A1(n3859), .A2(n3840), .ZN(n2226) );
  AND2_X1 U3135 ( .A1(n3), .A2(n113), .ZN(n2224) );
  AND2_X1 U3136 ( .A1(n3859), .A2(n113), .ZN(n2223) );
  OAI22_X1 U3137 ( .A1(n2171), .A2(n556), .B1(n2172), .B2(n559), .ZN(n3860) );
  NAND2_X1 U3138 ( .A1(n3858), .A2(n3837), .ZN(n2232) );
  NAND2_X1 U3139 ( .A1(n3859), .A2(n3837), .ZN(n2231) );
  AND2_X1 U3140 ( .A1(ADD_RS1[1]), .A2(n3861), .ZN(n3837) );
  NOR3_X1 U3141 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(ADD_RS1[0]), .ZN(n3859) );
  AND2_X1 U3142 ( .A1(n3841), .A2(n113), .ZN(n2229) );
  NOR2_X1 U3143 ( .A1(n3861), .A2(ADD_RS1[1]), .ZN(n3843) );
  INV_X1 U3144 ( .A(ADD_RS1[2]), .ZN(n3861) );
  NOR3_X1 U3145 ( .A1(n56), .A2(n84), .A3(n3844), .ZN(n3841) );
  INV_X1 U3146 ( .A(ADD_RS1[3]), .ZN(n3844) );
  AND2_X1 U3147 ( .A1(n3), .A2(n3838), .ZN(n2228) );
  NOR2_X1 U3148 ( .A1(ADD_RS1[1]), .A2(n57), .ZN(n3838) );
  NOR3_X1 U3149 ( .A1(ADD_RS1[3]), .A2(ADD_RS1[4]), .A3(n84), .ZN(n3858) );
  NAND2_X1 U3150 ( .A1(n3862), .A2(n437), .ZN(n2181) );
  AND3_X1 U3151 ( .A1(n715), .A2(ENABLE), .A3(RD1), .ZN(n2184) );
  INV_X1 U3152 ( .A(n3830), .ZN(n3862) );
  NAND4_X1 U3153 ( .A1(n3863), .A2(n3864), .A3(n3865), .A4(n3866), .ZN(n3830)
         );
  NOR3_X1 U3154 ( .A1(n3867), .A2(n1323), .A3(n3868), .ZN(n3866) );
  XNOR2_X1 U3155 ( .A(n1220), .B(ADD_RS1[1]), .ZN(n3868) );
  INV_X1 U3156 ( .A(ADD_WR[1]), .ZN(n1220) );
  OAI21_X1 U3157 ( .B1(n3869), .B2(n3870), .A(WR), .ZN(n1323) );
  NAND2_X1 U3158 ( .A1(n873), .A2(n874), .ZN(n3870) );
  INV_X1 U3159 ( .A(ADD_WR[4]), .ZN(n874) );
  INV_X1 U3160 ( .A(ADD_WR[3]), .ZN(n873) );
  INV_X1 U3161 ( .A(n910), .ZN(n3869) );
  NOR3_X1 U3162 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n910) );
  XNOR2_X1 U3163 ( .A(ADD_RS1[0]), .B(n1186), .ZN(n3867) );
  INV_X1 U3164 ( .A(ADD_WR[0]), .ZN(n1186) );
  XNOR2_X1 U3165 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n3865) );
  XNOR2_X1 U3166 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .ZN(n3864) );
  XNOR2_X1 U3167 ( .A(n57), .B(ADD_WR[2]), .ZN(n3863) );
endmodule


module Decode ( CLK, RST, Bubble, RF_WE, ZERO_FLAG, PC_IN, INS_IN, ADD_WR, 
        DATA_WR_IN, PC_OUT, A_OUT, B_OUT, IMM_OUT, ADD_RS1_HDU, ADD_RS2_HDU, 
        ADD_WR_OUT, ADD_RS1_OUT, ADD_RS2_OUT );
  input [31:0] PC_IN;
  input [31:0] INS_IN;
  input [4:0] ADD_WR;
  input [31:0] DATA_WR_IN;
  output [31:0] PC_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] ADD_RS1_HDU;
  output [4:0] ADD_RS2_HDU;
  output [4:0] ADD_WR_OUT;
  output [4:0] ADD_RS1_OUT;
  output [4:0] ADD_RS2_OUT;
  input CLK, RST, Bubble, RF_WE, ZERO_FLAG;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, sig_RST, sig_Rtype, sig_Itype,
         sig_Jtype, RD1, RD2, n6, n7, n11, n12;
  wire   [4:0] sig_ADD_WR;
  wire   [31:0] sig_IMM;
  wire   [4:0] sig_ADD_WRHAZ;
  wire   [4:0] sig_ADD_RS1HAZ;
  wire   [4:0] sig_ADD_RS2HAZ;

  NOR2_X2 U3 ( .A1(ZERO_FLAG), .A2(n12), .ZN(sig_RST) );
  instruction_type ins_type ( .INST_IN(INS_IN), .Rtype(sig_Rtype), .Itype(
        sig_Itype), .Jtype(sig_Jtype) );
  instruction_decomposition ins_dec ( .INST_IN({INS_IN[31], n7, n6, 
        INS_IN[28:0]}), .Rtype(sig_Rtype), .Itype(sig_Itype), .Jtype(sig_Jtype), .ADD_RS1({ADD_RS1_HDU[4], n13, n14, n15, ADD_RS1_HDU[0]}), .ADD_RS2({n16, 
        n17, n18, n19, n20}), .ADD_WR(sig_ADD_WR), .IMM(sig_IMM), .RD1(RD1), 
        .RD2(RD2) );
  regn_N32_7 regPC ( .DIN(PC_IN), .CLK(CLK), .EN(1'b1), .RST(sig_RST), .DOUT(
        PC_OUT) );
  regn_N32_6 regIMM ( .DIN(sig_IMM), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(IMM_OUT) );
  regn_N5_0 regWR ( .DIN(sig_ADD_WRHAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N5_4 regRS1 ( .DIN(sig_ADD_RS1HAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_RS1_OUT) );
  regn_N5_3 regRS2 ( .DIN(sig_ADD_RS2HAZ), .CLK(CLK), .EN(1'b1), .RST(sig_RST), 
        .DOUT(ADD_RS2_OUT) );
  mux21_NBIT5_0 muxRS1 ( .A(ADD_RS1_HDU), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .S(n11), .Z(sig_ADD_RS1HAZ) );
  mux21_NBIT5_2 muxRS2 ( .A(ADD_RS2_HDU), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .S(n11), .Z(sig_ADD_RS2HAZ) );
  mux21_NBIT5_1 muxWR ( .A(sig_ADD_WR), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .S(n11), .Z(sig_ADD_WRHAZ) );
  register_file_NBIT_ADD5_NBIT_DATA32 rf ( .CLK(CLK), .RST(RST), .ENABLE(1'b1), 
        .RD1(RD1), .RD2(RD2), .WR(RF_WE), .ADD_WR(ADD_WR), .ADD_RS1({
        ADD_RS1_HDU[4], n13, n14, n15, ADD_RS1_HDU[0]}), .ADD_RS2({n16, n17, 
        n18, n19, n20}), .DATAIN(DATA_WR_IN), .OUT1(A_OUT), .OUT2(B_OUT) );
  BUF_X1 U4 ( .A(Bubble), .Z(n11) );
  CLKBUF_X1 U5 ( .A(n18), .Z(ADD_RS2_HDU[2]) );
  CLKBUF_X1 U6 ( .A(n14), .Z(ADD_RS1_HDU[2]) );
  CLKBUF_X1 U7 ( .A(n19), .Z(ADD_RS2_HDU[1]) );
  CLKBUF_X1 U8 ( .A(n15), .Z(ADD_RS1_HDU[1]) );
  CLKBUF_X1 U9 ( .A(n20), .Z(ADD_RS2_HDU[0]) );
  CLKBUF_X1 U10 ( .A(INS_IN[29]), .Z(n6) );
  CLKBUF_X1 U11 ( .A(INS_IN[30]), .Z(n7) );
  CLKBUF_X1 U12 ( .A(n16), .Z(ADD_RS2_HDU[4]) );
  CLKBUF_X1 U13 ( .A(n17), .Z(ADD_RS2_HDU[3]) );
  CLKBUF_X1 U14 ( .A(n13), .Z(ADD_RS1_HDU[3]) );
  INV_X1 U15 ( .A(RST), .ZN(n12) );
endmodule


module Branch_Cond_Unit_NBIT32 ( RST, A, ALU_OPC, JUMP_TYPE, PC_SEL, ZERO );
  input [31:0] A;
  input [4:0] ALU_OPC;
  input [1:0] JUMP_TYPE;
  output [1:0] PC_SEL;
  input RST;
  output ZERO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n1, n2;

  NAND3_X1 U24 ( .A1(ALU_OPC[2]), .A2(n7), .A3(ALU_OPC[3]), .ZN(n9) );
  NAND3_X1 U25 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[2]), .A3(n20), .ZN(n7) );
  NOR4_X1 U3 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NOR4_X1 U4 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n19) );
  NOR4_X1 U5 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n14) );
  NOR4_X1 U6 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n18) );
  NOR4_X1 U7 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n13) );
  NOR4_X1 U8 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n17) );
  NOR4_X1 U9 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n12) );
  NOR2_X1 U10 ( .A1(n10), .A2(n11), .ZN(n8) );
  NAND4_X1 U11 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n10) );
  NAND4_X1 U12 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n11) );
  NOR4_X1 U13 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n16) );
  NOR3_X1 U14 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[4]), .A3(ALU_OPC[1]), .ZN(n20) );
  OAI211_X1 U15 ( .C1(n5), .C2(n6), .A(JUMP_TYPE[0]), .B(RST), .ZN(n4) );
  NOR2_X1 U16 ( .A1(n7), .A2(n1), .ZN(n6) );
  NOR4_X1 U17 ( .A1(n9), .A2(n8), .A3(ALU_OPC[4]), .A4(ALU_OPC[1]), .ZN(n5) );
  INV_X1 U18 ( .A(n8), .ZN(n1) );
  NAND2_X1 U19 ( .A1(JUMP_TYPE[1]), .A2(RST), .ZN(n3) );
  NAND2_X1 U20 ( .A1(n3), .A2(n4), .ZN(ZERO) );
  OAI22_X1 U21 ( .A1(JUMP_TYPE[0]), .A2(n3), .B1(JUMP_TYPE[1]), .B2(n4), .ZN(
        PC_SEL[0]) );
  NOR2_X1 U22 ( .A1(n2), .A2(n3), .ZN(PC_SEL[1]) );
  INV_X1 U23 ( .A(JUMP_TYPE[0]), .ZN(n2) );
endmodule


module ff_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module regn_N2 ( DIN, CLK, EN, RST, DOUT );
  input [1:0] DIN;
  output [1:0] DOUT;
  input CLK, EN, RST;
  wire   n1, n2, n3, n4, n5, n6;

  DFFR_X1 DOUT_reg_1_ ( .D(n6), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n4) );
  DFFR_X1 DOUT_reg_0_ ( .D(n5), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n3) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n4), .B2(EN), .A(n2), .ZN(n6) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
endmodule


module FWD_Unit ( RST, ADD_RS1, ADD_RS2, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, 
        RF_WE_WB, FWDA, FWDB );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  output [1:0] FWDA;
  output [1:0] FWDB;
  input RST, RF_WE_MEM, RF_WE_WB;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(FWDB[1]) );
  AOI21_X1 U4 ( .B1(n3), .B2(n4), .A(n5), .ZN(n1) );
  INV_X1 U5 ( .A(n6), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n2), .A2(n7), .ZN(FWDB[0]) );
  MUX2_X1 U7 ( .A(n6), .B(n8), .S(n5), .Z(n7) );
  AND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n5) );
  NOR2_X1 U9 ( .A1(n13), .A2(n14), .ZN(n12) );
  XOR2_X1 U10 ( .A(ADD_WR_MEM[4]), .B(ADD_RS2[4]), .Z(n14) );
  XOR2_X1 U11 ( .A(ADD_WR_MEM[3]), .B(ADD_RS2[3]), .Z(n13) );
  XNOR2_X1 U12 ( .A(ADD_RS2[1]), .B(ADD_WR_MEM[1]), .ZN(n11) );
  XNOR2_X1 U13 ( .A(ADD_RS2[2]), .B(ADD_WR_MEM[2]), .ZN(n10) );
  XNOR2_X1 U14 ( .A(ADD_RS2[0]), .B(ADD_WR_MEM[0]), .ZN(n9) );
  NAND4_X1 U15 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n6) );
  NOR2_X1 U16 ( .A1(n19), .A2(n20), .ZN(n18) );
  XOR2_X1 U17 ( .A(ADD_WR_WB[3]), .B(ADD_RS2[3]), .Z(n20) );
  XOR2_X1 U18 ( .A(ADD_WR_WB[2]), .B(ADD_RS2[2]), .Z(n19) );
  XNOR2_X1 U19 ( .A(ADD_RS2[4]), .B(ADD_WR_WB[4]), .ZN(n17) );
  XNOR2_X1 U20 ( .A(ADD_RS2[1]), .B(ADD_WR_WB[1]), .ZN(n16) );
  XNOR2_X1 U21 ( .A(ADD_RS2[0]), .B(ADD_WR_WB[0]), .ZN(n15) );
  NOR2_X1 U22 ( .A1(n21), .A2(n2), .ZN(FWDA[1]) );
  AOI21_X1 U23 ( .B1(n22), .B2(n4), .A(n23), .ZN(n21) );
  OAI21_X1 U24 ( .B1(n24), .B2(n25), .A(RF_WE_WB), .ZN(n4) );
  OR2_X1 U25 ( .A1(ADD_WR_WB[0]), .A2(ADD_WR_WB[1]), .ZN(n25) );
  OR3_X1 U26 ( .A1(ADD_WR_WB[3]), .A2(ADD_WR_WB[4]), .A3(ADD_WR_WB[2]), .ZN(
        n24) );
  INV_X1 U27 ( .A(n26), .ZN(n22) );
  NOR2_X1 U28 ( .A1(n2), .A2(n27), .ZN(FWDA[0]) );
  MUX2_X1 U29 ( .A(n26), .B(n8), .S(n23), .Z(n27) );
  AND4_X1 U30 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n23) );
  NOR2_X1 U31 ( .A1(n32), .A2(n33), .ZN(n31) );
  XOR2_X1 U32 ( .A(ADD_WR_MEM[4]), .B(ADD_RS1[4]), .Z(n33) );
  XOR2_X1 U33 ( .A(ADD_WR_MEM[3]), .B(ADD_RS1[3]), .Z(n32) );
  XNOR2_X1 U34 ( .A(ADD_RS1[1]), .B(ADD_WR_MEM[1]), .ZN(n30) );
  XNOR2_X1 U35 ( .A(ADD_RS1[2]), .B(ADD_WR_MEM[2]), .ZN(n29) );
  XNOR2_X1 U36 ( .A(ADD_RS1[0]), .B(ADD_WR_MEM[0]), .ZN(n28) );
  INV_X1 U37 ( .A(n34), .ZN(n8) );
  OAI21_X1 U38 ( .B1(n35), .B2(n36), .A(RF_WE_MEM), .ZN(n34) );
  OR2_X1 U39 ( .A1(ADD_WR_MEM[0]), .A2(ADD_WR_MEM[1]), .ZN(n36) );
  OR3_X1 U40 ( .A1(ADD_WR_MEM[3]), .A2(ADD_WR_MEM[4]), .A3(ADD_WR_MEM[2]), 
        .ZN(n35) );
  NAND4_X1 U41 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n26) );
  NOR2_X1 U42 ( .A1(n41), .A2(n42), .ZN(n40) );
  XOR2_X1 U43 ( .A(ADD_WR_WB[3]), .B(ADD_RS1[3]), .Z(n42) );
  XOR2_X1 U44 ( .A(ADD_WR_WB[2]), .B(ADD_RS1[2]), .Z(n41) );
  XNOR2_X1 U45 ( .A(ADD_RS1[4]), .B(ADD_WR_WB[4]), .ZN(n39) );
  XNOR2_X1 U46 ( .A(ADD_RS1[1]), .B(ADD_WR_WB[1]), .ZN(n38) );
  XNOR2_X1 U47 ( .A(ADD_RS1[0]), .B(ADD_WR_WB[0]), .ZN(n37) );
  INV_X1 U48 ( .A(RST), .ZN(n2) );
endmodule


module mux41_NBIT32_0 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  BUF_X1 U1 ( .A(n6), .Z(n72) );
  BUF_X1 U2 ( .A(n6), .Z(n73) );
  BUF_X1 U3 ( .A(n4), .Z(n78) );
  BUF_X1 U4 ( .A(n4), .Z(n79) );
  BUF_X1 U5 ( .A(n7), .Z(n1) );
  BUF_X1 U6 ( .A(n7), .Z(n70) );
  BUF_X1 U7 ( .A(n5), .Z(n75) );
  BUF_X1 U8 ( .A(n5), .Z(n76) );
  BUF_X1 U9 ( .A(n6), .Z(n74) );
  BUF_X1 U10 ( .A(n4), .Z(n80) );
  BUF_X1 U11 ( .A(n7), .Z(n71) );
  BUF_X1 U12 ( .A(n5), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n6) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n7) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n4) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n5) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n68), .A2(n69), .ZN(Z[0]) );
  AOI22_X1 U19 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n68) );
  AOI22_X1 U20 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n69) );
  NAND2_X1 U21 ( .A1(n44), .A2(n45), .ZN(Z[20]) );
  AOI22_X1 U22 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n44) );
  AOI22_X1 U23 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n45) );
  NAND2_X1 U24 ( .A1(n52), .A2(n53), .ZN(Z[17]) );
  AOI22_X1 U25 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n52) );
  AOI22_X1 U26 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n53) );
  NAND2_X1 U27 ( .A1(n60), .A2(n61), .ZN(Z[13]) );
  AOI22_X1 U28 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n60) );
  AOI22_X1 U29 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n61) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(Z[6]) );
  AOI22_X1 U31 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n12) );
  AOI22_X1 U32 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n13) );
  NAND2_X1 U33 ( .A1(n20), .A2(n21), .ZN(Z[31]) );
  AOI22_X1 U34 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n20) );
  AOI22_X1 U35 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n21) );
  NAND2_X1 U36 ( .A1(n28), .A2(n29), .ZN(Z[28]) );
  AOI22_X1 U37 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n28) );
  AOI22_X1 U38 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n29) );
  NAND2_X1 U39 ( .A1(n36), .A2(n37), .ZN(Z[24]) );
  AOI22_X1 U40 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n36) );
  AOI22_X1 U41 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n37) );
  NAND2_X1 U42 ( .A1(n42), .A2(n43), .ZN(Z[21]) );
  AOI22_X1 U43 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n42) );
  AOI22_X1 U44 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n43) );
  NAND2_X1 U45 ( .A1(n50), .A2(n51), .ZN(Z[18]) );
  AOI22_X1 U46 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n50) );
  AOI22_X1 U47 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n51) );
  NAND2_X1 U48 ( .A1(n58), .A2(n59), .ZN(Z[14]) );
  AOI22_X1 U49 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n58) );
  AOI22_X1 U50 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n59) );
  NAND2_X1 U51 ( .A1(n66), .A2(n67), .ZN(Z[10]) );
  AOI22_X1 U52 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n66) );
  AOI22_X1 U53 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n67) );
  NAND2_X1 U54 ( .A1(n10), .A2(n11), .ZN(Z[7]) );
  AOI22_X1 U55 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n10) );
  AOI22_X1 U56 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n11) );
  NAND2_X1 U57 ( .A1(n26), .A2(n27), .ZN(Z[29]) );
  AOI22_X1 U58 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n26) );
  AOI22_X1 U59 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n27) );
  NAND2_X1 U60 ( .A1(n34), .A2(n35), .ZN(Z[25]) );
  AOI22_X1 U61 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n34) );
  AOI22_X1 U62 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n35) );
  NAND2_X1 U63 ( .A1(n18), .A2(n19), .ZN(Z[3]) );
  AOI22_X1 U64 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n18) );
  AOI22_X1 U65 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n19) );
  NAND2_X1 U66 ( .A1(n40), .A2(n41), .ZN(Z[22]) );
  AOI22_X1 U67 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n40) );
  AOI22_X1 U68 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n41) );
  NAND2_X1 U69 ( .A1(n48), .A2(n49), .ZN(Z[19]) );
  AOI22_X1 U70 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n48) );
  AOI22_X1 U71 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n49) );
  NAND2_X1 U72 ( .A1(n56), .A2(n57), .ZN(Z[15]) );
  AOI22_X1 U73 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n56) );
  AOI22_X1 U74 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n57) );
  NAND2_X1 U75 ( .A1(n64), .A2(n65), .ZN(Z[11]) );
  AOI22_X1 U76 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n64) );
  AOI22_X1 U77 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n65) );
  NAND2_X1 U78 ( .A1(n8), .A2(n9), .ZN(Z[8]) );
  AOI22_X1 U79 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n8) );
  AOI22_X1 U80 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n9) );
  NAND2_X1 U81 ( .A1(n16), .A2(n17), .ZN(Z[4]) );
  AOI22_X1 U82 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n16) );
  AOI22_X1 U83 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n17) );
  NAND2_X1 U84 ( .A1(n24), .A2(n25), .ZN(Z[2]) );
  AOI22_X1 U85 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n24) );
  AOI22_X1 U86 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n25) );
  NAND2_X1 U87 ( .A1(n32), .A2(n33), .ZN(Z[26]) );
  AOI22_X1 U88 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n32) );
  AOI22_X1 U89 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n33) );
  NAND2_X1 U90 ( .A1(n38), .A2(n39), .ZN(Z[23]) );
  AOI22_X1 U91 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n38) );
  AOI22_X1 U92 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n39) );
  NAND2_X1 U93 ( .A1(n54), .A2(n55), .ZN(Z[16]) );
  AOI22_X1 U94 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n54) );
  AOI22_X1 U95 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n55) );
  NAND2_X1 U96 ( .A1(n62), .A2(n63), .ZN(Z[12]) );
  AOI22_X1 U97 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n62) );
  AOI22_X1 U98 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n63) );
  NAND2_X1 U99 ( .A1(n2), .A2(n3), .ZN(Z[9]) );
  AOI22_X1 U100 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n2) );
  AOI22_X1 U101 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n3) );
  NAND2_X1 U102 ( .A1(n14), .A2(n15), .ZN(Z[5]) );
  AOI22_X1 U103 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n14) );
  AOI22_X1 U104 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n15) );
  NAND2_X1 U105 ( .A1(n22), .A2(n23), .ZN(Z[30]) );
  AOI22_X1 U106 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n22) );
  AOI22_X1 U107 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n23) );
  NAND2_X1 U108 ( .A1(n30), .A2(n31), .ZN(Z[27]) );
  AOI22_X1 U109 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n30) );
  AOI22_X1 U110 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n31) );
  NAND2_X1 U111 ( .A1(n46), .A2(n47), .ZN(Z[1]) );
  AOI22_X1 U112 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n46) );
  AOI22_X1 U113 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n47) );
endmodule


module mux41_NBIT32_4 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n73) );
  BUF_X1 U2 ( .A(n147), .Z(n79) );
  BUF_X1 U3 ( .A(n144), .Z(n70) );
  BUF_X1 U4 ( .A(n146), .Z(n76) );
  BUF_X1 U5 ( .A(n145), .Z(n72) );
  BUF_X1 U6 ( .A(n147), .Z(n78) );
  BUF_X1 U7 ( .A(n144), .Z(n1) );
  BUF_X1 U8 ( .A(n146), .Z(n75) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NOR2_X1 U13 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U14 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U15 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U16 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U17 ( .A(S[0]), .ZN(n81) );
  NAND2_X1 U18 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  NAND2_X1 U19 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  NAND2_X1 U20 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  NAND2_X1 U21 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  AOI22_X1 U23 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  NAND2_X1 U24 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U25 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  AOI22_X1 U26 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  NAND2_X1 U27 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U28 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  AOI22_X1 U29 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  NAND2_X1 U30 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U31 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  AOI22_X1 U32 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  NAND2_X1 U33 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U34 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  AOI22_X1 U35 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  NAND2_X1 U36 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U37 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  AOI22_X1 U38 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  NAND2_X1 U39 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U40 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  AOI22_X1 U41 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  NAND2_X1 U42 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U43 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  AOI22_X1 U44 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  NAND2_X1 U45 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U46 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  AOI22_X1 U47 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  NAND2_X1 U48 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U49 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  AOI22_X1 U50 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  NAND2_X1 U51 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U52 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  AOI22_X1 U53 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  NAND2_X1 U54 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U55 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  AOI22_X1 U56 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  NAND2_X1 U57 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U58 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  AOI22_X1 U59 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  NAND2_X1 U60 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U61 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  AOI22_X1 U62 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  NAND2_X1 U63 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U64 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  AOI22_X1 U65 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  NAND2_X1 U66 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U67 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  AOI22_X1 U68 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  NAND2_X1 U69 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U70 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  AOI22_X1 U71 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  NAND2_X1 U72 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U73 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  AOI22_X1 U74 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  NAND2_X1 U75 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U76 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  AOI22_X1 U77 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  NAND2_X1 U78 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U79 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  AOI22_X1 U80 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  NAND2_X1 U81 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U82 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  AOI22_X1 U83 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  NAND2_X1 U84 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U85 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  AOI22_X1 U86 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  NAND2_X1 U87 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U88 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  AOI22_X1 U89 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  NAND2_X1 U90 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U91 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  AOI22_X1 U92 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  NAND2_X1 U93 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U94 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  AOI22_X1 U95 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  NAND2_X1 U96 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U97 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  AOI22_X1 U98 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  NAND2_X1 U99 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U100 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  AOI22_X1 U101 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  NAND2_X1 U102 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U103 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  AOI22_X1 U104 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  NAND2_X1 U105 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U106 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  AOI22_X1 U107 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U108 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  AOI22_X1 U109 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U110 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  AOI22_X1 U111 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U112 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U113 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
endmodule


module mux21_NBIT32_4 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U5 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U6 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U7 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U8 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U9 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U10 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U11 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U12 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U13 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U14 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U15 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U16 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U17 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U18 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U19 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U20 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U22 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U23 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U24 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U25 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U26 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U27 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U28 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U29 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U30 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U31 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U32 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U33 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U34 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U35 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U36 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U37 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U38 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U39 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U40 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U41 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U42 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U43 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U44 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U45 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U46 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U47 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U48 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U49 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U50 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U51 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U52 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U53 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U54 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U55 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U56 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U57 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U58 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U59 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U60 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U61 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U62 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U63 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U64 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U65 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module mux41_NBIT32_3 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n147), .Z(n78) );
  BUF_X1 U3 ( .A(n145), .Z(n73) );
  BUF_X1 U4 ( .A(n147), .Z(n79) );
  BUF_X1 U5 ( .A(n144), .Z(n1) );
  BUF_X1 U6 ( .A(n146), .Z(n75) );
  BUF_X1 U7 ( .A(n144), .Z(n70) );
  BUF_X1 U8 ( .A(n146), .Z(n76) );
  BUF_X1 U9 ( .A(n145), .Z(n74) );
  BUF_X1 U10 ( .A(n147), .Z(n80) );
  BUF_X1 U11 ( .A(n144), .Z(n71) );
  BUF_X1 U12 ( .A(n146), .Z(n77) );
  NAND2_X1 U13 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U14 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U15 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  NAND2_X1 U16 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U17 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  AOI22_X1 U18 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  NAND2_X1 U19 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  AOI22_X1 U21 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  NAND2_X1 U22 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U23 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  AOI22_X1 U24 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  NAND2_X1 U25 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U26 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  AOI22_X1 U27 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  NAND2_X1 U28 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U29 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  AOI22_X1 U30 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  NAND2_X1 U31 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U32 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  AOI22_X1 U33 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U35 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  AOI22_X1 U36 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  NAND2_X1 U37 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U38 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  AOI22_X1 U39 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  NAND2_X1 U40 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U41 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  AOI22_X1 U42 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  NAND2_X1 U43 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U44 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
  AOI22_X1 U45 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  NAND2_X1 U46 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U47 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  AOI22_X1 U48 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  NAND2_X1 U49 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U50 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  AOI22_X1 U51 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  NAND2_X1 U52 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U53 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  AOI22_X1 U54 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  NAND2_X1 U55 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U56 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  AOI22_X1 U57 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  NAND2_X1 U58 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U59 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  AOI22_X1 U60 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  NAND2_X1 U61 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U62 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  AOI22_X1 U63 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  NAND2_X1 U64 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U65 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  AOI22_X1 U66 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  NAND2_X1 U67 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U68 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  AOI22_X1 U69 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  NAND2_X1 U70 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U71 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  AOI22_X1 U72 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  NAND2_X1 U73 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U74 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  AOI22_X1 U75 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  NAND2_X1 U76 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U77 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  AOI22_X1 U78 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  NAND2_X1 U79 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U80 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  AOI22_X1 U81 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  NAND2_X1 U82 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U83 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  AOI22_X1 U84 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  NAND2_X1 U85 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U86 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  AOI22_X1 U87 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U88 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U89 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  AOI22_X1 U90 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  NAND2_X1 U91 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U92 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  AOI22_X1 U93 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  NAND2_X1 U94 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U95 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  AOI22_X1 U96 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  NAND2_X1 U97 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U98 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  AOI22_X1 U99 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  NAND2_X1 U100 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U101 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  AOI22_X1 U102 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  NAND2_X1 U103 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U104 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  AOI22_X1 U105 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  NAND2_X1 U106 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  AOI22_X1 U107 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  AOI22_X1 U108 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  NOR2_X1 U109 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  NOR2_X1 U110 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AND2_X1 U111 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  AND2_X1 U112 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  INV_X1 U113 ( .A(S[0]), .ZN(n81) );
endmodule


module comparator_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202;

  INV_X1 U1 ( .A(NE), .ZN(EQ) );
  INV_X1 U2 ( .A(n142), .ZN(n55) );
  INV_X1 U3 ( .A(n130), .ZN(n7) );
  INV_X1 U4 ( .A(n118), .ZN(n15) );
  INV_X1 U5 ( .A(n106), .ZN(n23) );
  INV_X1 U6 ( .A(n94), .ZN(n31) );
  INV_X1 U7 ( .A(n82), .ZN(n39) );
  INV_X1 U8 ( .A(n139), .ZN(n58) );
  INV_X1 U9 ( .A(n127), .ZN(n10) );
  INV_X1 U10 ( .A(n115), .ZN(n18) );
  INV_X1 U11 ( .A(n103), .ZN(n26) );
  INV_X1 U12 ( .A(n91), .ZN(n34) );
  INV_X1 U13 ( .A(n79), .ZN(n42) );
  INV_X1 U14 ( .A(GT), .ZN(LE) );
  INV_X1 U15 ( .A(n132), .ZN(n61) );
  INV_X1 U16 ( .A(n141), .ZN(n56) );
  INV_X1 U17 ( .A(n144), .ZN(n53) );
  INV_X1 U18 ( .A(n120), .ZN(n13) );
  INV_X1 U19 ( .A(n108), .ZN(n21) );
  INV_X1 U20 ( .A(n96), .ZN(n29) );
  INV_X1 U21 ( .A(n84), .ZN(n37) );
  INV_X1 U22 ( .A(n129), .ZN(n8) );
  INV_X1 U23 ( .A(n117), .ZN(n16) );
  INV_X1 U24 ( .A(n105), .ZN(n24) );
  INV_X1 U25 ( .A(n93), .ZN(n32) );
  INV_X1 U26 ( .A(n81), .ZN(n40) );
  INV_X1 U27 ( .A(n154), .ZN(n47) );
  INV_X1 U28 ( .A(n68), .ZN(n5) );
  INV_X1 U29 ( .A(A[30]), .ZN(n49) );
  INV_X1 U30 ( .A(n72), .ZN(n45) );
  INV_X1 U31 ( .A(n151), .ZN(n50) );
  INV_X1 U32 ( .A(B[30]), .ZN(n64) );
  INV_X1 U33 ( .A(n202), .ZN(n3) );
  INV_X1 U34 ( .A(B[1]), .ZN(n63) );
  INV_X1 U35 ( .A(A[0]), .ZN(n6) );
  INV_X1 U36 ( .A(A[3]), .ZN(n51) );
  INV_X1 U37 ( .A(A[5]), .ZN(n54) );
  INV_X1 U38 ( .A(A[7]), .ZN(n59) );
  INV_X1 U39 ( .A(A[9]), .ZN(n62) );
  INV_X1 U40 ( .A(A[11]), .ZN(n11) );
  INV_X1 U41 ( .A(A[13]), .ZN(n14) );
  INV_X1 U42 ( .A(A[15]), .ZN(n19) );
  INV_X1 U43 ( .A(B[31]), .ZN(n65) );
  INV_X1 U44 ( .A(A[17]), .ZN(n22) );
  INV_X1 U45 ( .A(A[19]), .ZN(n27) );
  INV_X1 U46 ( .A(A[21]), .ZN(n30) );
  INV_X1 U47 ( .A(A[23]), .ZN(n35) );
  INV_X1 U48 ( .A(A[25]), .ZN(n38) );
  INV_X1 U49 ( .A(A[27]), .ZN(n43) );
  INV_X1 U50 ( .A(A[29]), .ZN(n46) );
  INV_X1 U51 ( .A(A[4]), .ZN(n52) );
  INV_X1 U52 ( .A(A[8]), .ZN(n60) );
  INV_X1 U53 ( .A(A[12]), .ZN(n12) );
  INV_X1 U54 ( .A(A[2]), .ZN(n48) );
  INV_X1 U55 ( .A(A[6]), .ZN(n57) );
  INV_X1 U56 ( .A(A[10]), .ZN(n9) );
  INV_X1 U57 ( .A(A[14]), .ZN(n17) );
  INV_X1 U58 ( .A(A[16]), .ZN(n20) );
  INV_X1 U59 ( .A(A[20]), .ZN(n28) );
  INV_X1 U60 ( .A(A[24]), .ZN(n36) );
  INV_X1 U61 ( .A(A[28]), .ZN(n44) );
  INV_X1 U62 ( .A(A[18]), .ZN(n25) );
  INV_X1 U63 ( .A(A[22]), .ZN(n33) );
  INV_X1 U64 ( .A(A[26]), .ZN(n41) );
  INV_X1 U65 ( .A(GE), .ZN(LT) );
  NAND2_X1 U66 ( .A1(LE), .A2(GE), .ZN(NE) );
  AOI21_X1 U67 ( .B1(n66), .B2(n5), .A(n67), .ZN(GE) );
  AOI22_X1 U68 ( .A1(B[30]), .A2(n49), .B1(n69), .B2(n70), .ZN(n68) );
  AOI21_X1 U69 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U70 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U71 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U72 ( .B1(n80), .B2(n39), .A(n40), .ZN(n77) );
  AOI21_X1 U73 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U74 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U75 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U76 ( .B1(n92), .B2(n31), .A(n32), .ZN(n89) );
  AOI21_X1 U77 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U78 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U79 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U80 ( .B1(n104), .B2(n23), .A(n24), .ZN(n101) );
  AOI21_X1 U81 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U82 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U83 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U84 ( .B1(n116), .B2(n15), .A(n16), .ZN(n113) );
  AOI21_X1 U85 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U86 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U87 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U88 ( .B1(n128), .B2(n7), .A(n8), .ZN(n125) );
  AOI21_X1 U89 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U90 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U91 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U92 ( .B1(n140), .B2(n55), .A(n56), .ZN(n137) );
  AOI21_X1 U93 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U94 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U95 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U96 ( .B1(n152), .B2(n153), .A(n47), .ZN(n149) );
  AOI22_X1 U97 ( .A1(n155), .A2(n63), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U98 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U99 ( .A1(B[0]), .A2(n6), .ZN(n156) );
  OAI21_X1 U100 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  NAND2_X1 U101 ( .A1(A[31]), .A2(n65), .ZN(n66) );
  AOI22_X1 U102 ( .A1(A[30]), .A2(n64), .B1(n158), .B2(n70), .ZN(n157) );
  XOR2_X1 U103 ( .A(A[30]), .B(n64), .Z(n70) );
  AOI21_X1 U104 ( .B1(n159), .B2(n160), .A(n45), .ZN(n158) );
  NAND2_X1 U105 ( .A1(B[29]), .A2(n46), .ZN(n72) );
  OAI211_X1 U106 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NOR2_X1 U107 ( .A1(n163), .A2(n76), .ZN(n75) );
  AND2_X1 U108 ( .A1(B[28]), .A2(n44), .ZN(n76) );
  NAND2_X1 U109 ( .A1(B[27]), .A2(n43), .ZN(n78) );
  NAND2_X1 U110 ( .A1(n42), .A2(n164), .ZN(n162) );
  NOR2_X1 U111 ( .A1(n43), .A2(B[27]), .ZN(n79) );
  AOI211_X1 U112 ( .C1(n165), .C2(n166), .A(n82), .B(n37), .ZN(n161) );
  NAND2_X1 U113 ( .A1(B[25]), .A2(n38), .ZN(n84) );
  NAND2_X1 U114 ( .A1(n164), .A2(n81), .ZN(n82) );
  NAND2_X1 U115 ( .A1(B[26]), .A2(n41), .ZN(n81) );
  OR2_X1 U116 ( .A1(n41), .A2(B[26]), .ZN(n164) );
  OAI211_X1 U117 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NOR2_X1 U118 ( .A1(n169), .A2(n88), .ZN(n87) );
  AND2_X1 U119 ( .A1(B[24]), .A2(n36), .ZN(n88) );
  NAND2_X1 U120 ( .A1(B[23]), .A2(n35), .ZN(n90) );
  NAND2_X1 U121 ( .A1(n34), .A2(n170), .ZN(n168) );
  NOR2_X1 U122 ( .A1(n35), .A2(B[23]), .ZN(n91) );
  AOI211_X1 U123 ( .C1(n171), .C2(n172), .A(n94), .B(n29), .ZN(n167) );
  NAND2_X1 U124 ( .A1(B[21]), .A2(n30), .ZN(n96) );
  NAND2_X1 U125 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U126 ( .A1(B[22]), .A2(n33), .ZN(n93) );
  OR2_X1 U127 ( .A1(n33), .A2(B[22]), .ZN(n170) );
  OAI211_X1 U128 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NOR2_X1 U129 ( .A1(n175), .A2(n100), .ZN(n99) );
  AND2_X1 U130 ( .A1(B[20]), .A2(n28), .ZN(n100) );
  NAND2_X1 U131 ( .A1(B[19]), .A2(n27), .ZN(n102) );
  NAND2_X1 U132 ( .A1(n26), .A2(n176), .ZN(n174) );
  NOR2_X1 U133 ( .A1(n27), .A2(B[19]), .ZN(n103) );
  AOI211_X1 U134 ( .C1(n177), .C2(n178), .A(n106), .B(n21), .ZN(n173) );
  NAND2_X1 U135 ( .A1(B[17]), .A2(n22), .ZN(n108) );
  NAND2_X1 U136 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n25), .ZN(n105) );
  OR2_X1 U138 ( .A1(n25), .A2(B[18]), .ZN(n176) );
  OAI211_X1 U139 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NOR2_X1 U140 ( .A1(n181), .A2(n112), .ZN(n111) );
  AND2_X1 U141 ( .A1(B[16]), .A2(n20), .ZN(n112) );
  NAND2_X1 U142 ( .A1(B[15]), .A2(n19), .ZN(n114) );
  NAND2_X1 U143 ( .A1(n18), .A2(n182), .ZN(n180) );
  NOR2_X1 U144 ( .A1(n19), .A2(B[15]), .ZN(n115) );
  AOI211_X1 U145 ( .C1(n183), .C2(n184), .A(n118), .B(n13), .ZN(n179) );
  NAND2_X1 U146 ( .A1(B[13]), .A2(n14), .ZN(n120) );
  NAND2_X1 U147 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U148 ( .A1(B[14]), .A2(n17), .ZN(n117) );
  OR2_X1 U149 ( .A1(n17), .A2(B[14]), .ZN(n182) );
  OAI211_X1 U150 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NOR2_X1 U151 ( .A1(n187), .A2(n124), .ZN(n123) );
  AND2_X1 U152 ( .A1(B[12]), .A2(n12), .ZN(n124) );
  NAND2_X1 U153 ( .A1(B[11]), .A2(n11), .ZN(n126) );
  NAND2_X1 U154 ( .A1(n10), .A2(n188), .ZN(n186) );
  NOR2_X1 U155 ( .A1(n11), .A2(B[11]), .ZN(n127) );
  AOI211_X1 U156 ( .C1(n189), .C2(n190), .A(n130), .B(n61), .ZN(n185) );
  NAND2_X1 U157 ( .A1(B[9]), .A2(n62), .ZN(n132) );
  NAND2_X1 U158 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U159 ( .A1(B[10]), .A2(n9), .ZN(n129) );
  OR2_X1 U160 ( .A1(n9), .A2(B[10]), .ZN(n188) );
  OAI211_X1 U161 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NOR2_X1 U162 ( .A1(n193), .A2(n136), .ZN(n135) );
  AND2_X1 U163 ( .A1(B[8]), .A2(n60), .ZN(n136) );
  NAND2_X1 U164 ( .A1(B[7]), .A2(n59), .ZN(n138) );
  NAND2_X1 U165 ( .A1(n58), .A2(n194), .ZN(n192) );
  NOR2_X1 U166 ( .A1(n59), .A2(B[7]), .ZN(n139) );
  AOI211_X1 U167 ( .C1(n195), .C2(n196), .A(n142), .B(n53), .ZN(n191) );
  NAND2_X1 U168 ( .A1(B[5]), .A2(n54), .ZN(n144) );
  NAND2_X1 U169 ( .A1(n194), .A2(n141), .ZN(n142) );
  NAND2_X1 U170 ( .A1(B[6]), .A2(n57), .ZN(n141) );
  OR2_X1 U171 ( .A1(n57), .A2(B[6]), .ZN(n194) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NOR2_X1 U173 ( .A1(n198), .A2(n148), .ZN(n147) );
  AND2_X1 U174 ( .A1(B[4]), .A2(n52), .ZN(n148) );
  NAND2_X1 U175 ( .A1(B[3]), .A2(n51), .ZN(n150) );
  NAND3_X1 U176 ( .A1(n50), .A2(n199), .A3(n200), .ZN(n197) );
  OAI211_X1 U177 ( .C1(A[1]), .C2(n201), .A(n3), .B(n153), .ZN(n200) );
  AND2_X1 U178 ( .A1(n199), .A2(n154), .ZN(n153) );
  NAND2_X1 U179 ( .A1(B[2]), .A2(n48), .ZN(n154) );
  AOI21_X1 U180 ( .B1(A[1]), .B2(n201), .A(n63), .ZN(n202) );
  NOR2_X1 U181 ( .A1(n6), .A2(B[0]), .ZN(n201) );
  OR2_X1 U182 ( .A1(n48), .A2(B[2]), .ZN(n199) );
  NOR2_X1 U183 ( .A1(n51), .A2(B[3]), .ZN(n151) );
  NOR2_X1 U184 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U185 ( .A1(n54), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U186 ( .A1(n52), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U187 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U188 ( .A1(n62), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U189 ( .A1(n60), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U190 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U191 ( .A1(n14), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U192 ( .A1(n12), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U193 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U194 ( .A1(n22), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U195 ( .A1(n20), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U196 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U197 ( .A1(n30), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U198 ( .A1(n28), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U199 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U200 ( .A1(n38), .A2(B[25]), .ZN(n85) );
  NOR2_X1 U201 ( .A1(n36), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U202 ( .A1(n163), .A2(n73), .ZN(n159) );
  NOR2_X1 U203 ( .A1(n46), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U204 ( .A1(n44), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U205 ( .A1(n65), .A2(A[31]), .ZN(n67) );
endmodule


module comparator_NBIT32 ( A, B, OPSel, RES );
  input [31:0] A;
  input [31:0] B;
  input [2:0] OPSel;
  output [31:0] RES;
  wire   N26, N27, N28, N29, N30, N31, n15, n16, n17, n18, n19, n20, n2, n3,
         n4;
  assign RES[1] = 1'b0;
  assign RES[2] = 1'b0;
  assign RES[3] = 1'b0;
  assign RES[4] = 1'b0;
  assign RES[5] = 1'b0;
  assign RES[6] = 1'b0;
  assign RES[7] = 1'b0;
  assign RES[8] = 1'b0;
  assign RES[9] = 1'b0;
  assign RES[10] = 1'b0;
  assign RES[11] = 1'b0;
  assign RES[12] = 1'b0;
  assign RES[13] = 1'b0;
  assign RES[14] = 1'b0;
  assign RES[15] = 1'b0;
  assign RES[16] = 1'b0;
  assign RES[17] = 1'b0;
  assign RES[18] = 1'b0;
  assign RES[19] = 1'b0;
  assign RES[20] = 1'b0;
  assign RES[21] = 1'b0;
  assign RES[22] = 1'b0;
  assign RES[23] = 1'b0;
  assign RES[24] = 1'b0;
  assign RES[25] = 1'b0;
  assign RES[26] = 1'b0;
  assign RES[27] = 1'b0;
  assign RES[28] = 1'b0;
  assign RES[29] = 1'b0;
  assign RES[30] = 1'b0;
  assign RES[31] = 1'b0;

  comparator_NBIT32_DW01_cmp6_0 r57 ( .A(A), .B(B), .TC(1'b0), .LT(N30), .GT(
        N28), .EQ(N26), .LE(N31), .GE(N29), .NE(N27) );
  INV_X1 U3 ( .A(n15), .ZN(RES[0]) );
  AOI21_X1 U4 ( .B1(n16), .B2(n4), .A(n17), .ZN(n15) );
  INV_X1 U5 ( .A(OPSel[0]), .ZN(n3) );
  OAI22_X1 U6 ( .A1(n19), .A2(n2), .B1(OPSel[1]), .B2(n20), .ZN(n16) );
  INV_X1 U7 ( .A(OPSel[1]), .ZN(n2) );
  AOI22_X1 U8 ( .A1(N28), .A2(n3), .B1(N29), .B2(OPSel[0]), .ZN(n19) );
  AOI22_X1 U9 ( .A1(N26), .A2(n3), .B1(N27), .B2(OPSel[0]), .ZN(n20) );
  NOR3_X1 U10 ( .A1(n4), .A2(OPSel[1]), .A3(n18), .ZN(n17) );
  AOI22_X1 U11 ( .A1(N30), .A2(n3), .B1(OPSel[0]), .B2(N31), .ZN(n18) );
  INV_X1 U12 ( .A(OPSel[2]), .ZN(n4) );
endmodule


module shifter_NBIT32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input LOGIC_ARITH, LEFT_RIGHT;
  wire   n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n266, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649;

  AOI21_X2 U264 ( .B1(A[31]), .B2(B[18]), .A(n483), .ZN(n282) );
  OAI21_X2 U267 ( .B1(n613), .B2(n629), .A(n486), .ZN(n285) );
  AOI21_X2 U269 ( .B1(A[31]), .B2(n39), .A(n487), .ZN(n288) );
  AOI221_X2 U388 ( .B1(n31), .B2(A[18]), .C1(n21), .C2(A[17]), .A(n568), .ZN(
        n196) );
  NOR2_X2 U428 ( .A1(n639), .A2(n39), .ZN(n165) );
  NOR2_X2 U461 ( .A1(n643), .A2(n39), .ZN(n199) );
  NAND3_X1 U637 ( .A1(n227), .A2(n647), .A3(n228), .ZN(n226) );
  NAND3_X1 U638 ( .A1(n227), .A2(n647), .A3(B[4]), .ZN(n428) );
  NAND3_X1 U639 ( .A1(n445), .A2(n199), .A3(LEFT_RIGHT), .ZN(n240) );
  NAND3_X1 U641 ( .A1(n489), .A2(n629), .A3(n579), .ZN(n255) );
  NAND3_X1 U642 ( .A1(n267), .A2(n199), .A3(n445), .ZN(n138) );
  NOR4_X1 U2 ( .A1(B[20]), .A2(B[21]), .A3(B[19]), .A4(n594), .ZN(n484) );
  NOR2_X2 U3 ( .A1(n640), .A2(B[3]), .ZN(n262) );
  NOR2_X2 U4 ( .A1(n490), .A2(B[11]), .ZN(n283) );
  NAND3_X1 U5 ( .A1(n445), .A2(n35), .A3(LEFT_RIGHT), .ZN(n269) );
  INV_X1 U6 ( .A(n167), .ZN(n636) );
  NOR2_X1 U7 ( .A1(n637), .A2(B[4]), .ZN(n167) );
  INV_X1 U8 ( .A(n169), .ZN(n645) );
  INV_X1 U9 ( .A(n165), .ZN(n638) );
  INV_X1 U10 ( .A(n199), .ZN(n642) );
  INV_X1 U11 ( .A(n32), .ZN(n28) );
  INV_X1 U12 ( .A(n32), .ZN(n26) );
  INV_X1 U13 ( .A(n32), .ZN(n27) );
  INV_X1 U14 ( .A(n22), .ZN(n14) );
  INV_X1 U15 ( .A(n22), .ZN(n15) );
  INV_X1 U16 ( .A(n21), .ZN(n16) );
  INV_X1 U17 ( .A(n505), .ZN(n644) );
  INV_X1 U18 ( .A(n31), .ZN(n29) );
  INV_X1 U19 ( .A(n493), .ZN(n641) );
  NOR2_X1 U20 ( .A1(n646), .A2(n39), .ZN(n169) );
  NAND2_X1 U21 ( .A1(n488), .A2(n454), .ZN(n161) );
  INV_X1 U22 ( .A(n42), .ZN(n39) );
  OAI222_X1 U23 ( .A1(n79), .A2(n645), .B1(n63), .B2(n636), .C1(n91), .C2(n638), .ZN(n371) );
  OAI222_X1 U24 ( .A1(n82), .A2(n645), .B1(n62), .B2(n636), .C1(n95), .C2(n638), .ZN(n360) );
  OAI222_X1 U25 ( .A1(n85), .A2(n645), .B1(n73), .B2(n636), .C1(n99), .C2(n638), .ZN(n349) );
  OAI222_X1 U26 ( .A1(n87), .A2(n645), .B1(n76), .B2(n636), .C1(n104), .C2(
        n638), .ZN(n338) );
  NOR2_X1 U27 ( .A1(n41), .A2(n643), .ZN(n493) );
  OAI22_X1 U28 ( .A1(n116), .A2(n643), .B1(n127), .B2(n639), .ZN(n383) );
  INV_X1 U29 ( .A(n454), .ZN(n637) );
  AOI21_X1 U30 ( .B1(n135), .B2(n2), .A(n519), .ZN(n286) );
  AOI21_X1 U31 ( .B1(n130), .B2(n3), .A(n519), .ZN(n312) );
  BUF_X1 U32 ( .A(n138), .Z(n34) );
  BUF_X1 U33 ( .A(n138), .Z(n33) );
  NOR2_X1 U34 ( .A1(n383), .A2(n359), .ZN(n197) );
  NOR2_X1 U35 ( .A1(n119), .A2(n359), .ZN(n181) );
  BUF_X1 U36 ( .A(n138), .Z(n35) );
  NAND2_X1 U37 ( .A1(n488), .A2(n5), .ZN(n505) );
  INV_X1 U38 ( .A(n182), .ZN(n119) );
  INV_X1 U39 ( .A(n238), .ZN(n107) );
  INV_X1 U40 ( .A(n214), .ZN(n56) );
  INV_X1 U41 ( .A(n202), .ZN(n50) );
  INV_X1 U42 ( .A(n188), .ZN(n48) );
  NOR2_X1 U43 ( .A1(n613), .A2(n148), .ZN(n150) );
  OAI21_X2 U44 ( .B1(n612), .B2(n633), .A(n481), .ZN(n279) );
  NOR2_X1 U45 ( .A1(n640), .A2(n647), .ZN(n454) );
  NAND2_X1 U46 ( .A1(n484), .A2(n631), .ZN(n281) );
  AOI222_X1 U47 ( .A1(n370), .A2(n262), .B1(n320), .B2(n260), .C1(n185), .C2(
        n3), .ZN(n238) );
  INV_X1 U48 ( .A(n356), .ZN(n643) );
  AOI222_X1 U49 ( .A1(n168), .A2(n262), .B1(n355), .B2(n260), .C1(n170), .C2(
        n3), .ZN(n471) );
  AOI222_X1 U50 ( .A1(n402), .A2(n262), .B1(n403), .B2(n260), .C1(n464), .C2(
        n2), .ZN(n461) );
  NAND2_X1 U51 ( .A1(n488), .A2(n262), .ZN(n157) );
  NAND2_X1 U52 ( .A1(n488), .A2(n260), .ZN(n158) );
  OAI222_X1 U53 ( .A1(n374), .A2(n639), .B1(n646), .B2(n375), .C1(n376), .C2(
        n643), .ZN(n172) );
  OAI222_X1 U54 ( .A1(n132), .A2(n639), .B1(n362), .B2(n646), .C1(n363), .C2(
        n643), .ZN(n139) );
  OAI222_X1 U55 ( .A1(n614), .A2(n639), .B1(n293), .B2(n646), .C1(n405), .C2(
        n643), .ZN(n348) );
  OAI222_X1 U56 ( .A1(n616), .A2(n639), .B1(n46), .B2(n646), .C1(n387), .C2(
        n643), .ZN(n337) );
  AOI221_X1 U57 ( .B1(n130), .B2(n262), .C1(n355), .C2(n2), .A(n359), .ZN(n159) );
  AOI221_X1 U58 ( .B1(n135), .B2(n262), .C1(n403), .C2(n3), .A(n359), .ZN(n347) );
  OAI221_X1 U59 ( .B1(n106), .B2(n639), .C1(n90), .C2(n643), .A(n607), .ZN(
        n480) );
  AOI22_X1 U60 ( .A1(n454), .A2(n320), .B1(n260), .B2(n370), .ZN(n607) );
  AOI222_X1 U61 ( .A1(n169), .A2(n185), .B1(n493), .B2(n320), .C1(n167), .C2(
        n370), .ZN(n550) );
  OAI222_X1 U62 ( .A1(n62), .A2(n645), .B1(n363), .B2(n636), .C1(n82), .C2(
        n638), .ZN(n418) );
  OAI222_X1 U63 ( .A1(n73), .A2(n645), .B1(n405), .B2(n636), .C1(n85), .C2(
        n638), .ZN(n404) );
  OAI222_X1 U64 ( .A1(n76), .A2(n645), .B1(n387), .B2(n636), .C1(n87), .C2(
        n638), .ZN(n386) );
  INV_X1 U65 ( .A(n260), .ZN(n646) );
  NOR2_X1 U66 ( .A1(n648), .A2(B[4]), .ZN(n488) );
  INV_X1 U67 ( .A(n262), .ZN(n639) );
  INV_X1 U68 ( .A(n332), .ZN(n628) );
  OAI222_X1 U69 ( .A1(n133), .A2(n14), .B1(n29), .B2(n615), .C1(n1), .C2(n103), 
        .ZN(n602) );
  OAI221_X1 U70 ( .B1(n363), .B2(n639), .C1(n62), .C2(n643), .A(n522), .ZN(
        n314) );
  AOI22_X1 U71 ( .A1(n454), .A2(n58), .B1(n260), .B2(n420), .ZN(n522) );
  OAI221_X1 U72 ( .B1(n405), .B2(n639), .C1(n73), .C2(n643), .A(n509), .ZN(
        n290) );
  AOI22_X1 U73 ( .A1(n454), .A2(n52), .B1(n260), .B2(n407), .ZN(n509) );
  OAI221_X1 U74 ( .B1(n387), .B2(n639), .C1(n76), .C2(n643), .A(n496), .ZN(
        n271) );
  AOI22_X1 U75 ( .A1(n454), .A2(n390), .B1(n260), .B2(n389), .ZN(n496) );
  OAI21_X1 U76 ( .B1(n613), .B2(n631), .A(n486), .ZN(n253) );
  NOR2_X1 U77 ( .A1(n613), .A2(n647), .ZN(n359) );
  NOR2_X1 U78 ( .A1(n613), .A2(n2), .ZN(n519) );
  AOI221_X1 U79 ( .B1(n219), .B2(n199), .C1(n223), .C2(n39), .A(n224), .ZN(
        n222) );
  OAI222_X1 U80 ( .A1(n638), .A2(n71), .B1(n636), .B2(n93), .C1(n645), .C2(n81), .ZN(n224) );
  AOI221_X1 U81 ( .B1(n207), .B2(n199), .C1(n211), .C2(n39), .A(n212), .ZN(
        n210) );
  OAI222_X1 U82 ( .A1(n638), .A2(n68), .B1(n636), .B2(n97), .C1(n645), .C2(n84), .ZN(n212) );
  AOI221_X1 U83 ( .B1(n193), .B2(n199), .C1(n115), .C2(n39), .A(n200), .ZN(
        n198) );
  OAI222_X1 U84 ( .A1(n638), .A2(n75), .B1(n636), .B2(n101), .C1(n645), .C2(
        n196), .ZN(n200) );
  OAI22_X1 U85 ( .A1(n8), .A2(n131), .B1(n1), .B2(n266), .ZN(n533) );
  OAI221_X1 U86 ( .B1(n618), .B2(n642), .C1(n238), .C2(n41), .A(n239), .ZN(
        n229) );
  AOI222_X1 U87 ( .A1(n165), .A2(n178), .B1(n167), .B2(n186), .C1(n169), .C2(
        n184), .ZN(n239) );
  OAI221_X1 U88 ( .B1(n65), .B2(n642), .C1(n182), .C2(n41), .A(n183), .ZN(n173) );
  AOI222_X1 U89 ( .A1(n165), .A2(n184), .B1(n167), .B2(n185), .C1(n169), .C2(
        n186), .ZN(n183) );
  OAI221_X1 U90 ( .B1(n71), .B2(n642), .C1(n163), .C2(n42), .A(n164), .ZN(n141) );
  AOI222_X1 U91 ( .A1(n165), .A2(n166), .B1(n167), .B2(n168), .C1(n169), .C2(
        n170), .ZN(n164) );
  OAI221_X1 U92 ( .B1(n68), .B2(n642), .C1(n344), .C2(n42), .A(n581), .ZN(n572) );
  AOI222_X1 U93 ( .A1(n165), .A2(n516), .B1(n167), .B2(n402), .C1(n169), .C2(
        n464), .ZN(n581) );
  OAI221_X1 U94 ( .B1(n93), .B2(n638), .C1(n81), .C2(n642), .A(n534), .ZN(n526) );
  AOI222_X1 U95 ( .A1(n169), .A2(n168), .B1(n493), .B2(n129), .C1(n167), .C2(
        n355), .ZN(n534) );
  OAI221_X1 U96 ( .B1(n97), .B2(n638), .C1(n84), .C2(n642), .A(n520), .ZN(n511) );
  AOI222_X1 U97 ( .A1(n169), .A2(n402), .B1(n493), .B2(n134), .C1(n167), .C2(
        n403), .ZN(n520) );
  OAI221_X1 U98 ( .B1(n101), .B2(n638), .C1(n196), .C2(n642), .A(n507), .ZN(
        n498) );
  AOI222_X1 U99 ( .A1(n169), .A2(n453), .B1(n493), .B2(n382), .C1(n167), .C2(
        n506), .ZN(n507) );
  NOR2_X1 U100 ( .A1(n613), .A2(n8), .ZN(n382) );
  OAI221_X1 U101 ( .B1(n127), .B2(n161), .C1(n116), .C2(n158), .A(n162), .ZN(
        n503) );
  OAI221_X1 U102 ( .B1(n237), .B2(n160), .C1(n90), .C2(n161), .A(n162), .ZN(
        n235) );
  OAI221_X1 U103 ( .B1(n110), .B2(n160), .C1(n93), .C2(n161), .A(n162), .ZN(
        n220) );
  OAI221_X1 U104 ( .B1(n113), .B2(n160), .C1(n97), .C2(n161), .A(n162), .ZN(
        n208) );
  OAI221_X1 U105 ( .B1(n197), .B2(n160), .C1(n101), .C2(n161), .A(n162), .ZN(
        n194) );
  OAI221_X1 U106 ( .B1(n181), .B2(n160), .C1(n106), .C2(n161), .A(n162), .ZN(
        n179) );
  OAI221_X1 U107 ( .B1(n159), .B2(n160), .C1(n109), .C2(n161), .A(n162), .ZN(
        n155) );
  OAI221_X1 U108 ( .B1(n347), .B2(n160), .C1(n112), .C2(n161), .A(n162), .ZN(
        n577) );
  OAI221_X1 U109 ( .B1(n336), .B2(n160), .C1(n116), .C2(n161), .A(n162), .ZN(
        n560) );
  OAI221_X1 U110 ( .B1(n323), .B2(n160), .C1(n118), .C2(n161), .A(n162), .ZN(
        n548) );
  INV_X1 U111 ( .A(n370), .ZN(n118) );
  OAI221_X1 U112 ( .B1(n312), .B2(n160), .C1(n121), .C2(n161), .A(n162), .ZN(
        n531) );
  INV_X1 U113 ( .A(n355), .ZN(n121) );
  OAI221_X1 U114 ( .B1(n286), .B2(n160), .C1(n124), .C2(n161), .A(n162), .ZN(
        n517) );
  INV_X1 U115 ( .A(n403), .ZN(n124) );
  AND2_X1 U116 ( .A1(n491), .A2(n633), .ZN(n276) );
  AOI22_X1 U117 ( .A1(n480), .A2(n39), .B1(n43), .B2(n64), .ZN(n587) );
  INV_X1 U118 ( .A(n601), .ZN(n64) );
  AOI221_X1 U119 ( .B1(n4), .B2(n602), .C1(n454), .C2(n184), .A(n603), .ZN(
        n601) );
  OAI22_X1 U120 ( .A1(n618), .A2(n639), .B1(n65), .B2(n646), .ZN(n603) );
  AOI22_X1 U121 ( .A1(n420), .A2(n2), .B1(n58), .B2(n262), .ZN(n214) );
  AOI22_X1 U122 ( .A1(n407), .A2(n5), .B1(n52), .B2(n262), .ZN(n202) );
  AOI22_X1 U123 ( .A1(n389), .A2(n3), .B1(n390), .B2(n262), .ZN(n188) );
  AOI22_X1 U124 ( .A1(n168), .A2(n3), .B1(n355), .B2(n262), .ZN(n413) );
  AOI22_X1 U125 ( .A1(n402), .A2(n5), .B1(n403), .B2(n262), .ZN(n396) );
  AOI22_X1 U126 ( .A1(n452), .A2(n4), .B1(n453), .B2(n262), .ZN(n449) );
  AOI22_X1 U127 ( .A1(n370), .A2(n4), .B1(n320), .B2(n262), .ZN(n182) );
  AOI22_X1 U128 ( .A1(n355), .A2(n2), .B1(n129), .B2(n262), .ZN(n163) );
  AOI22_X1 U129 ( .A1(n403), .A2(n4), .B1(n134), .B2(n262), .ZN(n344) );
  AOI21_X1 U130 ( .B1(n148), .B2(n232), .A(n150), .ZN(n231) );
  OAI21_X1 U131 ( .B1(n233), .B2(n152), .A(n153), .ZN(n232) );
  AOI211_X1 U132 ( .C1(n644), .C2(n234), .A(n235), .B(n236), .ZN(n233) );
  OAI22_X1 U133 ( .A1(n65), .A2(n157), .B1(n78), .B2(n158), .ZN(n236) );
  AOI21_X1 U134 ( .B1(n148), .B2(n217), .A(n150), .ZN(n216) );
  OAI21_X1 U135 ( .B1(n218), .B2(n152), .A(n153), .ZN(n217) );
  AOI211_X1 U136 ( .C1(n644), .C2(n219), .A(n220), .B(n221), .ZN(n218) );
  OAI22_X1 U137 ( .A1(n71), .A2(n157), .B1(n81), .B2(n158), .ZN(n221) );
  AOI21_X1 U138 ( .B1(n148), .B2(n205), .A(n150), .ZN(n204) );
  OAI21_X1 U139 ( .B1(n206), .B2(n152), .A(n153), .ZN(n205) );
  AOI211_X1 U140 ( .C1(n644), .C2(n207), .A(n208), .B(n209), .ZN(n206) );
  OAI22_X1 U141 ( .A1(n68), .A2(n157), .B1(n84), .B2(n158), .ZN(n209) );
  AOI21_X1 U142 ( .B1(n148), .B2(n191), .A(n150), .ZN(n190) );
  OAI21_X1 U143 ( .B1(n192), .B2(n152), .A(n153), .ZN(n191) );
  AOI211_X1 U144 ( .C1(n644), .C2(n193), .A(n194), .B(n195), .ZN(n192) );
  OAI22_X1 U145 ( .A1(n75), .A2(n157), .B1(n196), .B2(n158), .ZN(n195) );
  AOI21_X1 U146 ( .B1(n148), .B2(n176), .A(n150), .ZN(n175) );
  OAI21_X1 U147 ( .B1(n177), .B2(n152), .A(n153), .ZN(n176) );
  AOI211_X1 U148 ( .C1(n644), .C2(n178), .A(n179), .B(n180), .ZN(n177) );
  OAI22_X1 U149 ( .A1(n78), .A2(n157), .B1(n90), .B2(n158), .ZN(n180) );
  AOI21_X1 U150 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  OAI21_X1 U151 ( .B1(n151), .B2(n152), .A(n153), .ZN(n149) );
  AOI211_X1 U152 ( .C1(n644), .C2(n154), .A(n155), .B(n156), .ZN(n151) );
  OAI22_X1 U153 ( .A1(n81), .A2(n157), .B1(n93), .B2(n158), .ZN(n156) );
  AOI21_X1 U154 ( .B1(n148), .B2(n575), .A(n150), .ZN(n574) );
  OAI21_X1 U155 ( .B1(n576), .B2(n152), .A(n153), .ZN(n575) );
  AOI211_X1 U156 ( .C1(n644), .C2(n305), .A(n577), .B(n578), .ZN(n576) );
  OAI22_X1 U157 ( .A1(n84), .A2(n157), .B1(n97), .B2(n158), .ZN(n578) );
  AOI21_X1 U158 ( .B1(n148), .B2(n558), .A(n150), .ZN(n557) );
  OAI21_X1 U159 ( .B1(n559), .B2(n152), .A(n153), .ZN(n558) );
  AOI211_X1 U160 ( .C1(n644), .C2(n261), .A(n560), .B(n561), .ZN(n559) );
  OAI22_X1 U161 ( .A1(n196), .A2(n157), .B1(n101), .B2(n158), .ZN(n561) );
  AOI21_X1 U162 ( .B1(n148), .B2(n546), .A(n150), .ZN(n545) );
  OAI21_X1 U163 ( .B1(n547), .B2(n152), .A(n153), .ZN(n546) );
  AOI211_X1 U164 ( .C1(n644), .C2(n184), .A(n548), .B(n549), .ZN(n547) );
  OAI22_X1 U165 ( .A1(n90), .A2(n157), .B1(n106), .B2(n158), .ZN(n549) );
  AOI21_X1 U166 ( .B1(n148), .B2(n529), .A(n150), .ZN(n528) );
  OAI21_X1 U167 ( .B1(n530), .B2(n152), .A(n153), .ZN(n529) );
  AOI211_X1 U168 ( .C1(n644), .C2(n166), .A(n531), .B(n532), .ZN(n530) );
  OAI22_X1 U169 ( .A1(n93), .A2(n157), .B1(n109), .B2(n158), .ZN(n532) );
  AOI21_X1 U170 ( .B1(n148), .B2(n514), .A(n150), .ZN(n513) );
  OAI21_X1 U171 ( .B1(n515), .B2(n152), .A(n153), .ZN(n514) );
  AOI211_X1 U172 ( .C1(n644), .C2(n516), .A(n517), .B(n518), .ZN(n515) );
  OAI22_X1 U173 ( .A1(n97), .A2(n157), .B1(n112), .B2(n158), .ZN(n518) );
  AOI21_X1 U174 ( .B1(n283), .B2(n415), .A(n285), .ZN(n414) );
  OAI21_X1 U175 ( .B1(n110), .B2(n287), .A(n288), .ZN(n415) );
  AOI21_X1 U176 ( .B1(n283), .B2(n398), .A(n285), .ZN(n397) );
  OAI21_X1 U177 ( .B1(n113), .B2(n287), .A(n288), .ZN(n398) );
  AOI21_X1 U178 ( .B1(n283), .B2(n385), .A(n285), .ZN(n384) );
  OAI21_X1 U179 ( .B1(n197), .B2(n287), .A(n288), .ZN(n385) );
  AOI21_X1 U180 ( .B1(n283), .B2(n369), .A(n285), .ZN(n368) );
  OAI21_X1 U181 ( .B1(n181), .B2(n287), .A(n288), .ZN(n369) );
  AOI21_X1 U182 ( .B1(n283), .B2(n335), .A(n285), .ZN(n334) );
  OAI21_X1 U183 ( .B1(n336), .B2(n287), .A(n288), .ZN(n335) );
  OAI211_X1 U184 ( .C1(n127), .C2(n646), .A(n401), .B(n449), .ZN(n257) );
  AOI21_X1 U185 ( .B1(n320), .B2(n4), .A(n519), .ZN(n323) );
  AOI21_X1 U186 ( .B1(n506), .B2(n5), .A(n519), .ZN(n336) );
  NAND2_X1 U187 ( .A1(n484), .A2(n633), .ZN(n249) );
  OAI21_X1 U188 ( .B1(n417), .B2(n637), .A(n471), .ZN(n440) );
  OAI21_X1 U189 ( .B1(n400), .B2(n637), .A(n461), .ZN(n302) );
  NOR2_X1 U190 ( .A1(n613), .A2(n484), .ZN(n483) );
  OAI21_X1 U191 ( .B1(n412), .B2(n637), .A(n471), .ZN(n434) );
  OAI21_X1 U192 ( .B1(n395), .B2(n637), .A(n461), .ZN(n297) );
  OAI21_X1 U193 ( .B1(n412), .B2(n646), .A(n413), .ZN(n223) );
  OAI21_X1 U194 ( .B1(n395), .B2(n646), .A(n396), .ZN(n211) );
  OAI21_X1 U195 ( .B1(n333), .B2(n647), .A(n449), .ZN(n246) );
  OAI21_X1 U196 ( .B1(n482), .B2(n281), .A(n282), .ZN(n479) );
  AOI21_X1 U197 ( .B1(n283), .B2(n485), .A(n285), .ZN(n482) );
  OAI21_X1 U198 ( .B1(n89), .B2(n287), .A(n288), .ZN(n485) );
  INV_X1 U199 ( .A(n480), .ZN(n89) );
  OAI21_X1 U200 ( .B1(n472), .B2(n281), .A(n282), .ZN(n470) );
  AOI21_X1 U201 ( .B1(n283), .B2(n473), .A(n285), .ZN(n472) );
  OAI21_X1 U202 ( .B1(n94), .B2(n287), .A(n288), .ZN(n473) );
  INV_X1 U203 ( .A(n440), .ZN(n94) );
  OAI21_X1 U204 ( .B1(n462), .B2(n281), .A(n282), .ZN(n460) );
  AOI21_X1 U205 ( .B1(n283), .B2(n463), .A(n285), .ZN(n462) );
  OAI21_X1 U206 ( .B1(n98), .B2(n287), .A(n288), .ZN(n463) );
  INV_X1 U207 ( .A(n302), .ZN(n98) );
  OAI21_X1 U208 ( .B1(n450), .B2(n281), .A(n282), .ZN(n448) );
  AOI21_X1 U209 ( .B1(n283), .B2(n451), .A(n285), .ZN(n450) );
  OAI21_X1 U210 ( .B1(n102), .B2(n287), .A(n288), .ZN(n451) );
  INV_X1 U211 ( .A(n257), .ZN(n102) );
  OAI21_X1 U212 ( .B1(n425), .B2(n281), .A(n282), .ZN(n424) );
  AOI21_X1 U213 ( .B1(n283), .B2(n426), .A(n285), .ZN(n425) );
  OAI21_X1 U214 ( .B1(n237), .B2(n287), .A(n288), .ZN(n426) );
  OAI21_X1 U215 ( .B1(n357), .B2(n281), .A(n282), .ZN(n354) );
  AOI21_X1 U216 ( .B1(n283), .B2(n358), .A(n285), .ZN(n357) );
  OAI21_X1 U217 ( .B1(n159), .B2(n287), .A(n288), .ZN(n358) );
  OAI21_X1 U218 ( .B1(n345), .B2(n281), .A(n282), .ZN(n343) );
  AOI21_X1 U219 ( .B1(n283), .B2(n346), .A(n285), .ZN(n345) );
  OAI21_X1 U220 ( .B1(n347), .B2(n287), .A(n288), .ZN(n346) );
  OAI21_X1 U221 ( .B1(n321), .B2(n281), .A(n282), .ZN(n319) );
  AOI21_X1 U222 ( .B1(n283), .B2(n322), .A(n285), .ZN(n321) );
  OAI21_X1 U223 ( .B1(n323), .B2(n287), .A(n288), .ZN(n322) );
  OAI21_X1 U224 ( .B1(n310), .B2(n281), .A(n282), .ZN(n309) );
  AOI21_X1 U225 ( .B1(n283), .B2(n311), .A(n285), .ZN(n310) );
  OAI21_X1 U226 ( .B1(n312), .B2(n287), .A(n288), .ZN(n311) );
  OAI21_X1 U227 ( .B1(n280), .B2(n281), .A(n282), .ZN(n277) );
  AOI21_X1 U228 ( .B1(n283), .B2(n284), .A(n285), .ZN(n280) );
  OAI21_X1 U229 ( .B1(n286), .B2(n287), .A(n288), .ZN(n284) );
  AOI22_X1 U230 ( .A1(n246), .A2(n39), .B1(n43), .B2(n247), .ZN(n245) );
  AOI22_X1 U231 ( .A1(n434), .A2(n39), .B1(n42), .B2(n435), .ZN(n433) );
  AOI22_X1 U232 ( .A1(n297), .A2(n39), .B1(n42), .B2(n298), .ZN(n296) );
  INV_X1 U233 ( .A(n452), .ZN(n101) );
  INV_X1 U234 ( .A(n464), .ZN(n97) );
  INV_X1 U235 ( .A(n170), .ZN(n93) );
  INV_X1 U236 ( .A(n186), .ZN(n90) );
  INV_X1 U237 ( .A(n516), .ZN(n84) );
  INV_X1 U238 ( .A(n166), .ZN(n81) );
  NOR2_X1 U239 ( .A1(n266), .A2(n8), .ZN(n580) );
  AOI21_X1 U240 ( .B1(n251), .B2(n438), .A(n253), .ZN(n437) );
  OAI21_X1 U241 ( .B1(n439), .B2(n255), .A(n256), .ZN(n438) );
  AOI22_X1 U242 ( .A1(n435), .A2(n40), .B1(B[4]), .B2(n440), .ZN(n439) );
  AOI21_X1 U243 ( .B1(n251), .B2(n300), .A(n253), .ZN(n299) );
  OAI21_X1 U244 ( .B1(n301), .B2(n255), .A(n256), .ZN(n300) );
  AOI22_X1 U245 ( .A1(n298), .A2(n40), .B1(B[4]), .B2(n302), .ZN(n301) );
  AOI21_X1 U246 ( .B1(n251), .B2(n252), .A(n253), .ZN(n248) );
  OAI21_X1 U247 ( .B1(n254), .B2(n255), .A(n256), .ZN(n252) );
  AOI22_X1 U248 ( .A1(n247), .A2(n40), .B1(B[4]), .B2(n257), .ZN(n254) );
  BUF_X1 U249 ( .A(n356), .Z(n2) );
  BUF_X1 U250 ( .A(n356), .Z(n3) );
  INV_X1 U251 ( .A(n293), .ZN(n52) );
  INV_X1 U252 ( .A(n184), .ZN(n78) );
  INV_X1 U253 ( .A(n506), .ZN(n127) );
  INV_X1 U254 ( .A(n185), .ZN(n106) );
  INV_X1 U255 ( .A(n412), .ZN(n129) );
  INV_X1 U256 ( .A(n395), .ZN(n134) );
  INV_X1 U257 ( .A(n390), .ZN(n46) );
  BUF_X1 U258 ( .A(n356), .Z(n4) );
  BUF_X1 U259 ( .A(n356), .Z(n5) );
  INV_X1 U260 ( .A(n453), .ZN(n116) );
  INV_X1 U261 ( .A(n154), .ZN(n71) );
  INV_X1 U262 ( .A(n305), .ZN(n68) );
  INV_X1 U263 ( .A(n178), .ZN(n65) );
  INV_X1 U265 ( .A(n168), .ZN(n109) );
  INV_X1 U266 ( .A(n402), .ZN(n112) );
  INV_X1 U268 ( .A(n261), .ZN(n75) );
  INV_X1 U270 ( .A(n419), .ZN(n82) );
  INV_X1 U271 ( .A(n406), .ZN(n85) );
  INV_X1 U272 ( .A(n388), .ZN(n87) );
  BUF_X1 U273 ( .A(n44), .Z(n42) );
  INV_X1 U274 ( .A(n362), .ZN(n58) );
  INV_X1 U275 ( .A(n474), .ZN(n62) );
  INV_X1 U276 ( .A(n465), .ZN(n73) );
  INV_X1 U277 ( .A(n455), .ZN(n76) );
  INV_X1 U278 ( .A(n267), .ZN(n8) );
  BUF_X1 U279 ( .A(n44), .Z(n43) );
  BUF_X1 U280 ( .A(n44), .Z(n40) );
  INV_X1 U281 ( .A(n417), .ZN(n130) );
  INV_X1 U282 ( .A(n400), .ZN(n135) );
  BUF_X1 U283 ( .A(n44), .Z(n41) );
  INV_X1 U284 ( .A(n373), .ZN(n79) );
  INV_X1 U285 ( .A(n420), .ZN(n132) );
  INV_X1 U286 ( .A(n407), .ZN(n614) );
  INV_X1 U287 ( .A(n389), .ZN(n616) );
  INV_X1 U288 ( .A(n429), .ZN(n63) );
  INV_X1 U289 ( .A(n372), .ZN(n91) );
  INV_X1 U290 ( .A(n361), .ZN(n95) );
  INV_X1 U291 ( .A(n350), .ZN(n99) );
  INV_X1 U292 ( .A(n339), .ZN(n104) );
  AND2_X1 U293 ( .A1(n238), .A2(n401), .ZN(n237) );
  INV_X1 U294 ( .A(n234), .ZN(n618) );
  INV_X1 U295 ( .A(n416), .ZN(n110) );
  OAI211_X1 U296 ( .C1(n417), .C2(n646), .A(n401), .B(n413), .ZN(n416) );
  INV_X1 U297 ( .A(n399), .ZN(n113) );
  OAI211_X1 U298 ( .C1(n400), .C2(n646), .A(n401), .B(n396), .ZN(n399) );
  INV_X1 U299 ( .A(n381), .ZN(n115) );
  AOI21_X1 U300 ( .B1(n260), .B2(n382), .A(n383), .ZN(n381) );
  OR4_X1 U301 ( .A1(B[21]), .A2(B[20]), .A3(B[19]), .A4(B[18]), .ZN(n598) );
  OAI22_X1 U302 ( .A1(n88), .A2(n1), .B1(n86), .B2(n8), .ZN(n568) );
  AOI222_X1 U303 ( .A1(n11), .A2(A[1]), .B1(A[0]), .B2(n18), .C1(n7), .C2(A[2]), .ZN(n293) );
  AOI221_X1 U304 ( .B1(n31), .B2(A[6]), .C1(n20), .C2(A[7]), .A(n525), .ZN(
        n363) );
  OAI22_X1 U305 ( .A1(n623), .A2(n1), .B1(n624), .B2(n8), .ZN(n525) );
  AOI221_X1 U306 ( .B1(n30), .B2(A[7]), .C1(n20), .C2(A[8]), .A(n570), .ZN(
        n405) );
  OAI22_X1 U307 ( .A1(n624), .A2(n1), .B1(n66), .B2(n8), .ZN(n570) );
  AOI221_X1 U308 ( .B1(n31), .B2(A[8]), .C1(n21), .C2(A[9]), .A(n552), .ZN(
        n387) );
  OAI22_X1 U309 ( .A1(n66), .A2(n1), .B1(n74), .B2(n8), .ZN(n552) );
  AOI221_X1 U310 ( .B1(n30), .B2(A[5]), .C1(n20), .C2(A[6]), .A(n541), .ZN(
        n376) );
  OAI22_X1 U311 ( .A1(n622), .A2(n1), .B1(n623), .B2(n8), .ZN(n541) );
  OAI221_X1 U312 ( .B1(n29), .B2(n613), .C1(n17), .C2(n266), .A(n609), .ZN(
        n320) );
  AOI22_X1 U313 ( .A1(A[29]), .A2(n10), .B1(A[28]), .B2(n267), .ZN(n609) );
  OAI221_X1 U314 ( .B1(n27), .B2(n128), .C1(n15), .C2(n126), .A(n535), .ZN(
        n355) );
  AOI22_X1 U315 ( .A1(A[26]), .A2(n11), .B1(A[25]), .B2(n6), .ZN(n535) );
  OAI221_X1 U316 ( .B1(n28), .B2(n131), .C1(n16), .C2(n128), .A(n585), .ZN(
        n403) );
  AOI22_X1 U317 ( .A1(A[27]), .A2(n9), .B1(A[26]), .B2(n267), .ZN(n585) );
  OR3_X1 U318 ( .A1(B[22]), .A2(B[24]), .A3(B[23]), .ZN(n594) );
  NAND3_X1 U319 ( .A1(n489), .A2(n629), .A3(n600), .ZN(n152) );
  NOR3_X1 U320 ( .A1(B[12]), .A2(B[14]), .A3(B[13]), .ZN(n600) );
  NAND3_X1 U321 ( .A1(n592), .A2(n632), .A3(n599), .ZN(n146) );
  INV_X1 U322 ( .A(B[22]), .ZN(n632) );
  NOR3_X1 U323 ( .A1(B[23]), .A2(B[25]), .A3(B[24]), .ZN(n599) );
  NAND2_X1 U324 ( .A1(A[31]), .A2(n648), .ZN(n162) );
  OAI221_X1 U325 ( .B1(n29), .B2(n86), .C1(n17), .C2(n83), .A(n606), .ZN(n184)
         );
  AOI22_X1 U326 ( .A1(A[13]), .A2(n10), .B1(A[12]), .B2(n267), .ZN(n606) );
  OAI221_X1 U327 ( .B1(n29), .B2(n126), .C1(n17), .C2(n123), .A(n608), .ZN(
        n370) );
  AOI22_X1 U328 ( .A1(A[25]), .A2(n10), .B1(A[24]), .B2(n267), .ZN(n608) );
  NAND2_X1 U329 ( .A1(n488), .A2(n489), .ZN(n287) );
  OAI221_X1 U330 ( .B1(n27), .B2(n117), .C1(n15), .C2(n114), .A(n536), .ZN(
        n168) );
  AOI22_X1 U331 ( .A1(A[22]), .A2(n9), .B1(A[21]), .B2(n7), .ZN(n536) );
  OAI221_X1 U332 ( .B1(n28), .B2(n120), .C1(n16), .C2(n117), .A(n583), .ZN(
        n402) );
  AOI22_X1 U333 ( .A1(A[23]), .A2(n9), .B1(A[22]), .B2(n267), .ZN(n583) );
  AOI221_X1 U334 ( .B1(A[1]), .B2(n32), .C1(A[2]), .C2(n18), .A(n540), .ZN(
        n374) );
  OAI22_X1 U335 ( .A1(n615), .A2(n1), .B1(n617), .B2(n8), .ZN(n540) );
  NAND2_X1 U336 ( .A1(A[31]), .A2(n152), .ZN(n153) );
  NAND2_X1 U337 ( .A1(A[31]), .A2(n146), .ZN(n147) );
  NOR2_X2 U338 ( .A1(n612), .A2(n591), .ZN(n144) );
  OAI221_X1 U339 ( .B1(n28), .B2(n266), .C1(n16), .C2(n131), .A(n564), .ZN(
        n506) );
  AOI22_X1 U340 ( .A1(A[28]), .A2(n9), .B1(A[27]), .B2(n7), .ZN(n564) );
  OAI221_X1 U341 ( .B1(n28), .B2(n123), .C1(n16), .C2(n120), .A(n565), .ZN(
        n453) );
  AOI22_X1 U342 ( .A1(A[24]), .A2(n9), .B1(A[23]), .B2(n7), .ZN(n565) );
  NOR2_X2 U343 ( .A1(n647), .A2(B[2]), .ZN(n260) );
  OAI221_X1 U344 ( .B1(n26), .B2(n114), .C1(n14), .C2(n111), .A(n611), .ZN(
        n185) );
  AOI22_X1 U345 ( .A1(A[21]), .A2(n11), .B1(A[20]), .B2(n6), .ZN(n611) );
  AOI222_X1 U346 ( .A1(n429), .A2(n5), .B1(n620), .B2(n262), .C1(n227), .C2(
        B[3]), .ZN(n327) );
  INV_X1 U347 ( .A(n376), .ZN(n620) );
  OAI221_X1 U348 ( .B1(n26), .B2(n77), .C1(n15), .C2(n74), .A(n444), .ZN(n154)
         );
  AOI22_X1 U349 ( .A1(A[10]), .A2(n11), .B1(A[9]), .B2(n6), .ZN(n444) );
  OAI221_X1 U350 ( .B1(n29), .B2(n80), .C1(n16), .C2(n77), .A(n586), .ZN(n305)
         );
  AOI22_X1 U351 ( .A1(A[11]), .A2(n10), .B1(A[10]), .B2(n267), .ZN(n586) );
  OAI221_X1 U352 ( .B1(n28), .B2(n83), .C1(n16), .C2(n80), .A(n567), .ZN(n261)
         );
  AOI22_X1 U353 ( .A1(A[12]), .A2(n9), .B1(A[11]), .B2(n7), .ZN(n567) );
  OAI221_X1 U354 ( .B1(n26), .B2(n623), .C1(n14), .C2(n622), .A(n443), .ZN(
        n219) );
  AOI22_X1 U355 ( .A1(A[6]), .A2(n11), .B1(A[5]), .B2(n7), .ZN(n443) );
  OAI221_X1 U356 ( .B1(n26), .B2(n624), .C1(n14), .C2(n623), .A(n306), .ZN(
        n207) );
  AOI22_X1 U357 ( .A1(A[7]), .A2(n11), .B1(A[6]), .B2(n6), .ZN(n306) );
  OAI221_X1 U358 ( .B1(n27), .B2(n66), .C1(n15), .C2(n624), .A(n265), .ZN(n193) );
  AOI22_X1 U359 ( .A1(A[8]), .A2(n10), .B1(A[7]), .B2(n6), .ZN(n265) );
  OAI221_X1 U360 ( .B1(n29), .B2(n100), .C1(n17), .C2(n96), .A(n610), .ZN(n186) );
  AOI22_X1 U361 ( .A1(A[17]), .A2(n10), .B1(A[16]), .B2(n267), .ZN(n610) );
  OAI221_X1 U362 ( .B1(n29), .B2(n74), .C1(n17), .C2(n66), .A(n604), .ZN(n178)
         );
  AOI22_X1 U363 ( .A1(A[9]), .A2(n10), .B1(A[8]), .B2(n267), .ZN(n604) );
  OAI221_X1 U364 ( .B1(n27), .B2(n88), .C1(n15), .C2(n86), .A(n537), .ZN(n166)
         );
  AOI22_X1 U365 ( .A1(A[14]), .A2(n11), .B1(A[13]), .B2(n7), .ZN(n537) );
  OAI221_X1 U366 ( .B1(n28), .B2(n92), .C1(n16), .C2(n88), .A(n584), .ZN(n516)
         );
  AOI22_X1 U367 ( .A1(A[15]), .A2(n9), .B1(A[14]), .B2(n7), .ZN(n584) );
  OAI221_X1 U368 ( .B1(n27), .B2(n80), .C1(n15), .C2(n83), .A(n494), .ZN(n373)
         );
  AOI22_X1 U369 ( .A1(A[15]), .A2(n9), .B1(A[16]), .B2(n6), .ZN(n494) );
  OAI221_X1 U370 ( .B1(n27), .B2(n133), .C1(n15), .C2(n615), .A(n523), .ZN(
        n420) );
  AOI22_X1 U371 ( .A1(A[4]), .A2(n10), .B1(A[5]), .B2(n7), .ZN(n523) );
  OAI221_X1 U372 ( .B1(n28), .B2(n615), .C1(n16), .C2(n617), .A(n571), .ZN(
        n407) );
  AOI22_X1 U373 ( .A1(A[5]), .A2(n9), .B1(A[6]), .B2(n7), .ZN(n571) );
  OAI221_X1 U374 ( .B1(n28), .B2(n617), .C1(n16), .C2(n619), .A(n554), .ZN(
        n389) );
  AOI22_X1 U375 ( .A1(A[6]), .A2(n9), .B1(A[7]), .B2(n7), .ZN(n554) );
  OAI221_X1 U376 ( .B1(n49), .B2(n29), .C1(n103), .C2(n14), .A(n553), .ZN(n390) );
  AOI22_X1 U377 ( .A1(A[2]), .A2(n9), .B1(A[3]), .B2(n7), .ZN(n553) );
  OAI221_X1 U378 ( .B1(n28), .B2(n624), .C1(n16), .C2(n66), .A(n542), .ZN(n429) );
  AOI22_X1 U379 ( .A1(A[11]), .A2(n9), .B1(A[12]), .B2(n7), .ZN(n542) );
  OAI221_X1 U380 ( .B1(n28), .B2(n111), .C1(n16), .C2(n108), .A(n566), .ZN(
        n452) );
  AOI22_X1 U381 ( .A1(A[20]), .A2(n9), .B1(A[19]), .B2(n7), .ZN(n566) );
  OAI221_X1 U382 ( .B1(n28), .B2(n105), .C1(n16), .C2(n100), .A(n538), .ZN(
        n170) );
  AOI22_X1 U383 ( .A1(A[18]), .A2(n9), .B1(A[17]), .B2(n7), .ZN(n538) );
  OAI221_X1 U384 ( .B1(n28), .B2(n108), .C1(n16), .C2(n105), .A(n582), .ZN(
        n464) );
  AOI22_X1 U385 ( .A1(A[19]), .A2(n10), .B1(A[18]), .B2(n7), .ZN(n582) );
  INV_X1 U386 ( .A(A[31]), .ZN(n613) );
  AOI22_X1 U387 ( .A1(n267), .A2(A[1]), .B1(n11), .B2(A[0]), .ZN(n362) );
  NAND2_X1 U389 ( .A1(B[4]), .A2(n579), .ZN(n160) );
  OAI222_X1 U390 ( .A1(n79), .A2(n636), .B1(n326), .B2(n642), .C1(n91), .C2(
        n645), .ZN(n325) );
  AOI222_X1 U391 ( .A1(A[27]), .A2(n10), .B1(A[25]), .B2(n30), .C1(A[26]), 
        .C2(n18), .ZN(n326) );
  AOI222_X1 U392 ( .A1(A[28]), .A2(n10), .B1(A[26]), .B2(n30), .C1(A[27]), 
        .C2(n19), .ZN(n316) );
  AOI222_X1 U393 ( .A1(A[29]), .A2(n11), .B1(A[27]), .B2(n32), .C1(A[28]), 
        .C2(n18), .ZN(n292) );
  AOI222_X1 U394 ( .A1(A[30]), .A2(n11), .B1(A[28]), .B2(n30), .C1(A[29]), 
        .C2(n22), .ZN(n273) );
  AOI21_X1 U395 ( .B1(A[31]), .B2(B[11]), .A(n487), .ZN(n256) );
  AOI21_X1 U396 ( .B1(A[31]), .B2(B[25]), .A(n483), .ZN(n250) );
  OAI222_X1 U397 ( .A1(n171), .A2(n36), .B1(n55), .B2(n626), .C1(n623), .C2(
        n33), .ZN(RES[8]) );
  INV_X1 U398 ( .A(n172), .ZN(n55) );
  AOI221_X1 U399 ( .B1(n140), .B2(n173), .C1(n142), .C2(n174), .A(n144), .ZN(
        n171) );
  OAI21_X1 U400 ( .B1(n175), .B2(n146), .A(n147), .ZN(n174) );
  OAI222_X1 U401 ( .A1(n187), .A2(n36), .B1(n188), .B2(n626), .C1(n622), .C2(
        n33), .ZN(RES[7]) );
  AOI221_X1 U402 ( .B1(n140), .B2(n61), .C1(n142), .C2(n189), .A(n144), .ZN(
        n187) );
  INV_X1 U403 ( .A(n198), .ZN(n61) );
  OAI21_X1 U404 ( .B1(n190), .B2(n146), .A(n147), .ZN(n189) );
  OAI222_X1 U405 ( .A1(n136), .A2(n36), .B1(n59), .B2(n626), .C1(n624), .C2(
        n33), .ZN(RES[9]) );
  INV_X1 U406 ( .A(n139), .ZN(n59) );
  AOI221_X1 U407 ( .B1(n140), .B2(n141), .C1(n142), .C2(n143), .A(n144), .ZN(
        n136) );
  OAI21_X1 U408 ( .B1(n145), .B2(n146), .A(n147), .ZN(n143) );
  OAI222_X1 U409 ( .A1(n539), .A2(n36), .B1(n327), .B2(n626), .C1(n77), .C2(
        n35), .ZN(RES[12]) );
  AOI221_X1 U410 ( .B1(n140), .B2(n543), .C1(n142), .C2(n544), .A(n144), .ZN(
        n539) );
  OAI21_X1 U411 ( .B1(n545), .B2(n146), .A(n147), .ZN(n544) );
  OAI221_X1 U412 ( .B1(n90), .B2(n638), .C1(n78), .C2(n642), .A(n550), .ZN(
        n543) );
  OAI222_X1 U413 ( .A1(n521), .A2(n36), .B1(n57), .B2(n626), .C1(n80), .C2(n35), .ZN(RES[13]) );
  INV_X1 U414 ( .A(n314), .ZN(n57) );
  AOI221_X1 U415 ( .B1(n140), .B2(n526), .C1(n142), .C2(n527), .A(n144), .ZN(
        n521) );
  OAI21_X1 U416 ( .B1(n528), .B2(n146), .A(n147), .ZN(n527) );
  OAI222_X1 U417 ( .A1(n508), .A2(n36), .B1(n51), .B2(n626), .C1(n83), .C2(n35), .ZN(RES[14]) );
  INV_X1 U418 ( .A(n290), .ZN(n51) );
  AOI221_X1 U419 ( .B1(n140), .B2(n511), .C1(n142), .C2(n512), .A(n144), .ZN(
        n508) );
  OAI21_X1 U420 ( .B1(n513), .B2(n146), .A(n147), .ZN(n512) );
  OAI222_X1 U421 ( .A1(n551), .A2(n36), .B1(n45), .B2(n626), .C1(n74), .C2(n35), .ZN(RES[11]) );
  INV_X1 U422 ( .A(n337), .ZN(n45) );
  AOI221_X1 U423 ( .B1(n140), .B2(n555), .C1(n142), .C2(n556), .A(n144), .ZN(
        n551) );
  OAI21_X1 U424 ( .B1(n557), .B2(n146), .A(n147), .ZN(n556) );
  OAI222_X1 U425 ( .A1(n495), .A2(n36), .B1(n47), .B2(n626), .C1(n86), .C2(n35), .ZN(RES[15]) );
  INV_X1 U426 ( .A(n271), .ZN(n47) );
  AOI221_X1 U427 ( .B1(n140), .B2(n498), .C1(n142), .C2(n499), .A(n144), .ZN(
        n495) );
  OAI21_X1 U429 ( .B1(n500), .B2(n146), .A(n147), .ZN(n499) );
  OAI222_X1 U430 ( .A1(n569), .A2(n36), .B1(n53), .B2(n626), .C1(n66), .C2(n35), .ZN(RES[10]) );
  INV_X1 U431 ( .A(n348), .ZN(n53) );
  AOI221_X1 U432 ( .B1(n140), .B2(n572), .C1(n142), .C2(n573), .A(n144), .ZN(
        n569) );
  OAI21_X1 U433 ( .B1(n574), .B2(n146), .A(n147), .ZN(n573) );
  OAI222_X1 U434 ( .A1(n201), .A2(n36), .B1(n202), .B2(n626), .C1(n621), .C2(
        n33), .ZN(RES[6]) );
  AOI221_X1 U435 ( .B1(n140), .B2(n67), .C1(n142), .C2(n203), .A(n144), .ZN(
        n201) );
  INV_X1 U436 ( .A(n210), .ZN(n67) );
  OAI21_X1 U437 ( .B1(n204), .B2(n146), .A(n147), .ZN(n203) );
  OAI222_X1 U438 ( .A1(n213), .A2(n36), .B1(n214), .B2(n626), .C1(n619), .C2(
        n33), .ZN(RES[5]) );
  AOI221_X1 U439 ( .B1(n140), .B2(n70), .C1(n142), .C2(n215), .A(n144), .ZN(
        n213) );
  INV_X1 U440 ( .A(n222), .ZN(n70) );
  OAI21_X1 U441 ( .B1(n216), .B2(n146), .A(n147), .ZN(n215) );
  OAI221_X1 U442 ( .B1(n27), .B2(n83), .C1(n15), .C2(n86), .A(n476), .ZN(n419)
         );
  AOI22_X1 U443 ( .A1(A[16]), .A2(n11), .B1(A[17]), .B2(n6), .ZN(n476) );
  OAI221_X1 U444 ( .B1(n27), .B2(n86), .C1(n15), .C2(n88), .A(n467), .ZN(n406)
         );
  AOI22_X1 U445 ( .A1(A[17]), .A2(n9), .B1(A[18]), .B2(n7), .ZN(n467) );
  OAI221_X1 U446 ( .B1(n27), .B2(n88), .C1(n15), .C2(n92), .A(n457), .ZN(n388)
         );
  AOI22_X1 U447 ( .A1(A[18]), .A2(n10), .B1(A[19]), .B2(n6), .ZN(n457) );
  OAI221_X1 U448 ( .B1(n26), .B2(n92), .C1(n14), .C2(n96), .A(n430), .ZN(n372)
         );
  AOI22_X1 U449 ( .A1(A[19]), .A2(n11), .B1(A[20]), .B2(n6), .ZN(n430) );
  OAI221_X1 U450 ( .B1(n29), .B2(n622), .C1(n17), .C2(n621), .A(n605), .ZN(
        n234) );
  AOI22_X1 U451 ( .A1(A[5]), .A2(n10), .B1(A[4]), .B2(n267), .ZN(n605) );
  OAI221_X1 U452 ( .B1(n258), .B2(n643), .C1(n196), .C2(n637), .A(n259), .ZN(
        n247) );
  AOI22_X1 U453 ( .A1(n260), .A2(n261), .B1(n262), .B2(n193), .ZN(n259) );
  AOI222_X1 U454 ( .A1(A[4]), .A2(n11), .B1(A[6]), .B2(n31), .C1(A[5]), .C2(
        n19), .ZN(n258) );
  OAI221_X1 U455 ( .B1(n303), .B2(n643), .C1(n84), .C2(n637), .A(n304), .ZN(
        n298) );
  AOI22_X1 U456 ( .A1(n260), .A2(n305), .B1(n262), .B2(n207), .ZN(n304) );
  AOI222_X1 U457 ( .A1(A[3]), .A2(n10), .B1(A[5]), .B2(n32), .C1(A[4]), .C2(
        n19), .ZN(n303) );
  OAI221_X1 U458 ( .B1(n441), .B2(n643), .C1(n81), .C2(n637), .A(n442), .ZN(
        n435) );
  AOI22_X1 U459 ( .A1(n260), .A2(n154), .B1(n262), .B2(n219), .ZN(n442) );
  AOI222_X1 U460 ( .A1(A[2]), .A2(n10), .B1(A[4]), .B2(n30), .C1(A[3]), .C2(
        n20), .ZN(n441) );
  INV_X1 U462 ( .A(n228), .ZN(n626) );
  OAI221_X1 U463 ( .B1(n27), .B2(n66), .C1(n15), .C2(n74), .A(n524), .ZN(n474)
         );
  AOI22_X1 U464 ( .A1(A[12]), .A2(n11), .B1(A[13]), .B2(n7), .ZN(n524) );
  OAI221_X1 U465 ( .B1(n27), .B2(n74), .C1(n15), .C2(n77), .A(n510), .ZN(n465)
         );
  AOI22_X1 U466 ( .A1(A[13]), .A2(n9), .B1(A[14]), .B2(n6), .ZN(n510) );
  OAI221_X1 U467 ( .B1(n27), .B2(n77), .C1(n15), .C2(n80), .A(n497), .ZN(n455)
         );
  AOI22_X1 U468 ( .A1(A[14]), .A2(n10), .B1(A[15]), .B2(n7), .ZN(n497) );
  OAI221_X1 U469 ( .B1(n26), .B2(n96), .C1(n14), .C2(n100), .A(n421), .ZN(n361) );
  AOI22_X1 U470 ( .A1(A[20]), .A2(n11), .B1(A[21]), .B2(n6), .ZN(n421) );
  OAI221_X1 U471 ( .B1(n26), .B2(n100), .C1(n14), .C2(n105), .A(n408), .ZN(
        n350) );
  AOI22_X1 U472 ( .A1(A[21]), .A2(n11), .B1(A[22]), .B2(n6), .ZN(n408) );
  OAI221_X1 U473 ( .B1(n26), .B2(n105), .C1(n14), .C2(n108), .A(n391), .ZN(
        n339) );
  AOI22_X1 U474 ( .A1(A[22]), .A2(n9), .B1(A[23]), .B2(n6), .ZN(n391) );
  OAI221_X1 U475 ( .B1(n26), .B2(n108), .C1(n14), .C2(n111), .A(n377), .ZN(
        n324) );
  AOI22_X1 U476 ( .A1(A[23]), .A2(n9), .B1(A[24]), .B2(n6), .ZN(n377) );
  OAI221_X1 U477 ( .B1(n26), .B2(n111), .C1(n14), .C2(n114), .A(n364), .ZN(
        n313) );
  AOI22_X1 U478 ( .A1(A[24]), .A2(n10), .B1(A[25]), .B2(n6), .ZN(n364) );
  OAI221_X1 U479 ( .B1(n26), .B2(n114), .C1(n14), .C2(n117), .A(n351), .ZN(
        n289) );
  AOI22_X1 U480 ( .A1(A[25]), .A2(n11), .B1(A[26]), .B2(n6), .ZN(n351) );
  OAI221_X1 U481 ( .B1(n26), .B2(n117), .C1(n14), .C2(n120), .A(n340), .ZN(
        n270) );
  AOI22_X1 U482 ( .A1(A[26]), .A2(n10), .B1(A[27]), .B2(n6), .ZN(n340) );
  AOI22_X1 U483 ( .A1(n640), .A2(n506), .B1(B[2]), .B2(n382), .ZN(n333) );
  AOI21_X1 U484 ( .B1(n22), .B2(A[31]), .A(n533), .ZN(n412) );
  AOI21_X1 U485 ( .B1(n11), .B2(A[31]), .A(n580), .ZN(n395) );
  AOI21_X1 U486 ( .B1(B[1]), .B2(A[31]), .A(n533), .ZN(n417) );
  AOI21_X1 U487 ( .B1(n8), .B2(A[31]), .A(n580), .ZN(n400) );
  NOR2_X1 U488 ( .A1(n490), .A2(B[18]), .ZN(n251) );
  OAI22_X1 U489 ( .A1(B[2]), .A2(n374), .B1(n640), .B2(n375), .ZN(n227) );
  OAI221_X1 U490 ( .B1(n196), .B2(n638), .C1(n75), .C2(n642), .A(n562), .ZN(
        n555) );
  AOI221_X1 U491 ( .B1(n169), .B2(n452), .C1(n167), .C2(n453), .A(n563), .ZN(
        n562) );
  NOR3_X1 U492 ( .A1(n41), .A2(B[3]), .A3(n333), .ZN(n563) );
  NOR2_X1 U493 ( .A1(B[0]), .A2(B[1]), .ZN(n267) );
  AOI21_X1 U494 ( .B1(n634), .B2(n590), .A(n144), .ZN(n481) );
  INV_X1 U495 ( .A(n592), .ZN(n634) );
  NAND2_X1 U496 ( .A1(A[31]), .A2(n490), .ZN(n486) );
  OAI221_X1 U497 ( .B1(n225), .B2(n36), .C1(n617), .C2(n33), .A(n226), .ZN(
        RES[4]) );
  AOI221_X1 U498 ( .B1(n140), .B2(n229), .C1(n142), .C2(n230), .A(n144), .ZN(
        n225) );
  OAI21_X1 U499 ( .B1(n231), .B2(n146), .A(n147), .ZN(n230) );
  NAND2_X1 U500 ( .A1(n454), .A2(A[31]), .ZN(n401) );
  NOR2_X1 U501 ( .A1(B[2]), .A2(B[3]), .ZN(n356) );
  AOI21_X1 U502 ( .B1(n148), .B2(n501), .A(n150), .ZN(n500) );
  OAI21_X1 U503 ( .B1(n502), .B2(n152), .A(n153), .ZN(n501) );
  AOI211_X1 U504 ( .C1(B[4]), .C2(A[31]), .A(n503), .B(n504), .ZN(n502) );
  OAI22_X1 U505 ( .A1(n196), .A2(n505), .B1(n101), .B2(n157), .ZN(n504) );
  INV_X1 U506 ( .A(A[10]), .ZN(n66) );
  OAI21_X1 U507 ( .B1(n489), .B2(n613), .A(n162), .ZN(n487) );
  NOR3_X1 U508 ( .A1(n332), .A2(B[3]), .A3(n333), .ZN(n331) );
  INV_X1 U509 ( .A(B[3]), .ZN(n647) );
  INV_X1 U510 ( .A(A[11]), .ZN(n74) );
  INV_X1 U511 ( .A(A[15]), .ZN(n86) );
  INV_X1 U512 ( .A(A[9]), .ZN(n624) );
  INV_X1 U513 ( .A(A[16]), .ZN(n88) );
  BUF_X1 U514 ( .A(n137), .Z(n36) );
  BUF_X1 U515 ( .A(n137), .Z(n37) );
  NAND2_X1 U516 ( .A1(A[0]), .A2(n6), .ZN(n375) );
  INV_X1 U517 ( .A(A[23]), .ZN(n114) );
  INV_X1 U518 ( .A(A[19]), .ZN(n100) );
  INV_X1 U519 ( .A(A[24]), .ZN(n117) );
  INV_X1 U520 ( .A(A[20]), .ZN(n105) );
  INV_X1 U521 ( .A(A[21]), .ZN(n108) );
  INV_X1 U522 ( .A(A[22]), .ZN(n111) );
  INV_X1 U523 ( .A(A[8]), .ZN(n623) );
  INV_X1 U524 ( .A(A[12]), .ZN(n77) );
  INV_X1 U525 ( .A(A[13]), .ZN(n80) );
  INV_X1 U526 ( .A(A[14]), .ZN(n83) );
  INV_X1 U527 ( .A(A[30]), .ZN(n266) );
  INV_X1 U528 ( .A(A[3]), .ZN(n615) );
  OR4_X1 U529 ( .A1(B[13]), .A2(B[14]), .A3(B[12]), .A4(n596), .ZN(n490) );
  OR3_X1 U530 ( .A1(B[15]), .A2(B[17]), .A3(B[16]), .ZN(n596) );
  INV_X1 U531 ( .A(B[2]), .ZN(n640) );
  INV_X1 U532 ( .A(A[17]), .ZN(n92) );
  INV_X1 U533 ( .A(A[7]), .ZN(n622) );
  INV_X1 U534 ( .A(A[18]), .ZN(n96) );
  INV_X1 U535 ( .A(A[25]), .ZN(n120) );
  AND3_X1 U536 ( .A1(n579), .A2(n591), .A3(n597), .ZN(n445) );
  NOR3_X1 U537 ( .A1(n152), .A2(n146), .A3(n630), .ZN(n597) );
  INV_X1 U538 ( .A(n148), .ZN(n630) );
  INV_X1 U539 ( .A(A[4]), .ZN(n617) );
  INV_X1 U540 ( .A(n590), .ZN(n612) );
  INV_X1 U541 ( .A(A[27]), .ZN(n126) );
  INV_X1 U542 ( .A(A[26]), .ZN(n123) );
  INV_X1 U543 ( .A(A[6]), .ZN(n621) );
  INV_X1 U544 ( .A(A[5]), .ZN(n619) );
  INV_X1 U545 ( .A(A[28]), .ZN(n128) );
  INV_X1 U546 ( .A(A[29]), .ZN(n131) );
  INV_X1 U547 ( .A(B[25]), .ZN(n633) );
  INV_X1 U548 ( .A(A[2]), .ZN(n133) );
  AND2_X1 U549 ( .A1(n140), .A2(n199), .ZN(n278) );
  INV_X1 U550 ( .A(A[1]), .ZN(n103) );
  INV_X1 U551 ( .A(n579), .ZN(n648) );
  INV_X1 U552 ( .A(A[0]), .ZN(n49) );
  OR2_X1 U553 ( .A1(n625), .A2(B[1]), .ZN(n1) );
  NAND2_X1 U554 ( .A1(n140), .A2(n40), .ZN(n332) );
  INV_X1 U555 ( .A(n436), .ZN(n627) );
  NAND2_X1 U556 ( .A1(B[1]), .A2(B[0]), .ZN(n263) );
  NAND2_X1 U557 ( .A1(B[1]), .A2(n625), .ZN(n264) );
  INV_X1 U558 ( .A(B[11]), .ZN(n629) );
  INV_X1 U559 ( .A(B[18]), .ZN(n631) );
  AND2_X1 U560 ( .A1(n142), .A2(n592), .ZN(n491) );
  BUF_X1 U561 ( .A(n137), .Z(n38) );
  INV_X1 U562 ( .A(B[0]), .ZN(n625) );
  INV_X1 U563 ( .A(B[4]), .ZN(n44) );
  NOR2_X2 U564 ( .A1(n635), .A2(LOGIC_ARITH), .ZN(n142) );
  INV_X1 U565 ( .A(n591), .ZN(n635) );
  NOR3_X1 U566 ( .A1(B[9]), .A2(B[8]), .A3(B[10]), .ZN(n489) );
  NOR3_X1 U567 ( .A1(B[7]), .A2(B[6]), .A3(B[5]), .ZN(n579) );
  NOR3_X1 U568 ( .A1(B[28]), .A2(B[27]), .A3(B[26]), .ZN(n592) );
  OAI222_X1 U569 ( .A1(n468), .A2(n269), .B1(n469), .B2(n37), .C1(n92), .C2(
        n34), .ZN(RES[17]) );
  AOI221_X1 U570 ( .B1(n165), .B2(n474), .C1(n199), .C2(n419), .A(n475), .ZN(
        n468) );
  AOI221_X1 U571 ( .B1(n276), .B2(n470), .C1(n628), .C2(n434), .A(n279), .ZN(
        n469) );
  OAI222_X1 U572 ( .A1(n132), .A2(n636), .B1(n362), .B2(n641), .C1(n363), .C2(
        n645), .ZN(n475) );
  OAI222_X1 U573 ( .A1(n458), .A2(n269), .B1(n459), .B2(n38), .C1(n96), .C2(
        n34), .ZN(RES[18]) );
  AOI221_X1 U574 ( .B1(n165), .B2(n465), .C1(n199), .C2(n406), .A(n466), .ZN(
        n458) );
  AOI221_X1 U575 ( .B1(n276), .B2(n460), .C1(n628), .C2(n297), .A(n279), .ZN(
        n459) );
  OAI222_X1 U576 ( .A1(n614), .A2(n636), .B1(n293), .B2(n641), .C1(n405), .C2(
        n645), .ZN(n466) );
  OAI222_X1 U577 ( .A1(n446), .A2(n269), .B1(n447), .B2(n37), .C1(n100), .C2(
        n34), .ZN(RES[19]) );
  AOI221_X1 U578 ( .B1(n165), .B2(n455), .C1(n199), .C2(n388), .A(n456), .ZN(
        n446) );
  AOI221_X1 U579 ( .B1(n276), .B2(n448), .C1(n628), .C2(n246), .A(n279), .ZN(
        n447) );
  OAI222_X1 U580 ( .A1(n616), .A2(n636), .B1(n46), .B2(n641), .C1(n387), .C2(
        n645), .ZN(n456) );
  OAI222_X1 U581 ( .A1(n422), .A2(n269), .B1(n423), .B2(n37), .C1(n105), .C2(
        n34), .ZN(RES[20]) );
  AOI221_X1 U582 ( .B1(n165), .B2(n373), .C1(n199), .C2(n372), .A(n427), .ZN(
        n422) );
  AOI221_X1 U583 ( .B1(n276), .B2(n424), .C1(n628), .C2(n107), .A(n279), .ZN(
        n423) );
  OAI221_X1 U584 ( .B1(n376), .B2(n636), .C1(n63), .C2(n645), .A(n428), .ZN(
        n427) );
  OAI222_X1 U585 ( .A1(n409), .A2(n269), .B1(n410), .B2(n37), .C1(n108), .C2(
        n34), .ZN(RES[21]) );
  AOI221_X1 U586 ( .B1(n276), .B2(n411), .C1(n628), .C2(n223), .A(n279), .ZN(
        n410) );
  AOI221_X1 U587 ( .B1(n199), .B2(n361), .C1(B[4]), .C2(n56), .A(n418), .ZN(
        n409) );
  OAI21_X1 U588 ( .B1(n414), .B2(n281), .A(n282), .ZN(n411) );
  OAI222_X1 U589 ( .A1(n392), .A2(n269), .B1(n393), .B2(n37), .C1(n111), .C2(
        n34), .ZN(RES[22]) );
  AOI221_X1 U590 ( .B1(n276), .B2(n394), .C1(n628), .C2(n211), .A(n279), .ZN(
        n393) );
  AOI221_X1 U591 ( .B1(n199), .B2(n350), .C1(B[4]), .C2(n50), .A(n404), .ZN(
        n392) );
  OAI21_X1 U592 ( .B1(n397), .B2(n281), .A(n282), .ZN(n394) );
  OAI222_X1 U593 ( .A1(n378), .A2(n269), .B1(n379), .B2(n37), .C1(n114), .C2(
        n34), .ZN(RES[23]) );
  AOI221_X1 U594 ( .B1(n276), .B2(n380), .C1(n628), .C2(n115), .A(n279), .ZN(
        n379) );
  AOI221_X1 U595 ( .B1(n199), .B2(n339), .C1(B[4]), .C2(n48), .A(n386), .ZN(
        n378) );
  OAI21_X1 U596 ( .B1(n384), .B2(n281), .A(n282), .ZN(n380) );
  OAI222_X1 U597 ( .A1(n365), .A2(n269), .B1(n366), .B2(n37), .C1(n117), .C2(
        n34), .ZN(RES[24]) );
  AOI221_X1 U598 ( .B1(n276), .B2(n367), .C1(n628), .C2(n119), .A(n279), .ZN(
        n366) );
  AOI221_X1 U599 ( .B1(n199), .B2(n324), .C1(n39), .C2(n172), .A(n371), .ZN(
        n365) );
  OAI21_X1 U600 ( .B1(n368), .B2(n281), .A(n282), .ZN(n367) );
  OAI222_X1 U601 ( .A1(n352), .A2(n269), .B1(n353), .B2(n37), .C1(n120), .C2(
        n34), .ZN(RES[25]) );
  AOI221_X1 U602 ( .B1(n276), .B2(n354), .C1(n628), .C2(n122), .A(n279), .ZN(
        n353) );
  AOI221_X1 U603 ( .B1(n199), .B2(n313), .C1(n39), .C2(n139), .A(n360), .ZN(
        n352) );
  INV_X1 U604 ( .A(n163), .ZN(n122) );
  OAI222_X1 U605 ( .A1(n477), .A2(n269), .B1(n478), .B2(n38), .C1(n88), .C2(
        n35), .ZN(RES[16]) );
  AOI221_X1 U606 ( .B1(n165), .B2(n429), .C1(n199), .C2(n373), .A(n492), .ZN(
        n477) );
  AOI221_X1 U607 ( .B1(n276), .B2(n479), .C1(n628), .C2(n480), .A(n279), .ZN(
        n478) );
  OAI222_X1 U608 ( .A1(n374), .A2(n636), .B1(n375), .B2(n641), .C1(n376), .C2(
        n645), .ZN(n492) );
  OAI222_X1 U609 ( .A1(n341), .A2(n269), .B1(n342), .B2(n37), .C1(n123), .C2(
        n34), .ZN(RES[26]) );
  AOI221_X1 U610 ( .B1(n276), .B2(n343), .C1(n628), .C2(n125), .A(n279), .ZN(
        n342) );
  AOI221_X1 U611 ( .B1(n199), .B2(n289), .C1(n39), .C2(n348), .A(n349), .ZN(
        n341) );
  INV_X1 U612 ( .A(n344), .ZN(n125) );
  OAI222_X1 U613 ( .A1(n328), .A2(n269), .B1(n329), .B2(n37), .C1(n126), .C2(
        n34), .ZN(RES[27]) );
  AOI211_X1 U614 ( .C1(n276), .C2(n330), .A(n279), .B(n331), .ZN(n329) );
  AOI221_X1 U615 ( .B1(n199), .B2(n270), .C1(n39), .C2(n337), .A(n338), .ZN(
        n328) );
  OAI21_X1 U616 ( .B1(n334), .B2(n281), .A(n282), .ZN(n330) );
  OAI222_X1 U617 ( .A1(n317), .A2(n269), .B1(n318), .B2(n37), .C1(n128), .C2(
        n34), .ZN(RES[28]) );
  AOI221_X1 U618 ( .B1(n165), .B2(n324), .C1(n39), .C2(n54), .A(n325), .ZN(
        n317) );
  AOI221_X1 U619 ( .B1(n276), .B2(n319), .C1(n278), .C2(n320), .A(n279), .ZN(
        n318) );
  INV_X1 U620 ( .A(n327), .ZN(n54) );
  OAI222_X1 U621 ( .A1(n307), .A2(n269), .B1(n308), .B2(n37), .C1(n131), .C2(
        n33), .ZN(RES[29]) );
  AOI221_X1 U622 ( .B1(n165), .B2(n313), .C1(n39), .C2(n314), .A(n315), .ZN(
        n307) );
  AOI221_X1 U623 ( .B1(n276), .B2(n309), .C1(n278), .C2(n129), .A(n279), .ZN(
        n308) );
  OAI222_X1 U624 ( .A1(n82), .A2(n636), .B1(n316), .B2(n642), .C1(n95), .C2(
        n645), .ZN(n315) );
  OAI222_X1 U625 ( .A1(n274), .A2(n269), .B1(n275), .B2(n38), .C1(n266), .C2(
        n33), .ZN(RES[30]) );
  AOI221_X1 U626 ( .B1(n165), .B2(n289), .C1(n39), .C2(n290), .A(n291), .ZN(
        n274) );
  AOI221_X1 U627 ( .B1(n276), .B2(n277), .C1(n278), .C2(n134), .A(n279), .ZN(
        n275) );
  OAI222_X1 U628 ( .A1(n85), .A2(n636), .B1(n292), .B2(n642), .C1(n99), .C2(
        n645), .ZN(n291) );
  OAI221_X1 U629 ( .B1(n293), .B2(n240), .C1(n133), .C2(n33), .A(n294), .ZN(
        RES[2]) );
  AOI221_X1 U630 ( .B1(n242), .B2(n295), .C1(n627), .C2(n69), .A(n244), .ZN(
        n294) );
  INV_X1 U631 ( .A(n296), .ZN(n69) );
  OAI21_X1 U632 ( .B1(n299), .B2(n249), .A(n250), .ZN(n295) );
  OAI221_X1 U633 ( .B1(n362), .B2(n240), .C1(n103), .C2(n33), .A(n431), .ZN(
        RES[1]) );
  AOI221_X1 U634 ( .B1(n242), .B2(n432), .C1(n627), .C2(n72), .A(n244), .ZN(
        n431) );
  INV_X1 U635 ( .A(n433), .ZN(n72) );
  OAI21_X1 U636 ( .B1(n437), .B2(n249), .A(n250), .ZN(n432) );
  OAI221_X1 U640 ( .B1(n46), .B2(n240), .C1(n615), .C2(n33), .A(n241), .ZN(
        RES[3]) );
  AOI221_X1 U643 ( .B1(n242), .B2(n243), .C1(n627), .C2(n60), .A(n244), .ZN(
        n241) );
  INV_X1 U644 ( .A(n245), .ZN(n60) );
  OAI21_X1 U645 ( .B1(n248), .B2(n249), .A(n250), .ZN(n243) );
  NOR2_X1 U646 ( .A1(B[29]), .A2(B[30]), .ZN(n591) );
  AND2_X1 U647 ( .A1(LOGIC_ARITH), .A2(n445), .ZN(n140) );
  NOR2_X1 U648 ( .A1(n613), .A2(LOGIC_ARITH), .ZN(n590) );
  OAI221_X1 U649 ( .B1(n587), .B2(n436), .C1(n49), .C2(n33), .A(n588), .ZN(
        RES[0]) );
  NOR2_X1 U650 ( .A1(n269), .A2(n39), .ZN(n228) );
  AOI21_X1 U651 ( .B1(n242), .B2(n589), .A(n244), .ZN(n588) );
  OAI21_X1 U652 ( .B1(n593), .B2(n249), .A(n250), .ZN(n589) );
  AOI21_X1 U653 ( .B1(n251), .B2(n595), .A(n253), .ZN(n593) );
  OAI21_X1 U654 ( .B1(n587), .B2(n255), .A(n256), .ZN(n595) );
  AND2_X1 U655 ( .A1(n491), .A2(n649), .ZN(n242) );
  NAND2_X1 U656 ( .A1(n35), .A2(n649), .ZN(n137) );
  NAND2_X1 U657 ( .A1(n140), .A2(n649), .ZN(n436) );
  NOR2_X1 U658 ( .A1(n481), .A2(LEFT_RIGHT), .ZN(n244) );
  INV_X1 U659 ( .A(LEFT_RIGHT), .ZN(n649) );
  OAI222_X1 U660 ( .A1(n268), .A2(n269), .B1(LEFT_RIGHT), .B2(n612), .C1(n613), 
        .C2(n34), .ZN(RES[31]) );
  AOI221_X1 U661 ( .B1(n165), .B2(n270), .C1(n39), .C2(n271), .A(n272), .ZN(
        n268) );
  OAI222_X1 U662 ( .A1(n87), .A2(n636), .B1(n273), .B2(n642), .C1(n104), .C2(
        n645), .ZN(n272) );
  NOR4_X4 U663 ( .A1(B[16]), .A2(B[17]), .A3(B[15]), .A4(n598), .ZN(n148) );
  INV_X1 U664 ( .A(n8), .ZN(n6) );
  INV_X1 U665 ( .A(n8), .ZN(n7) );
  INV_X1 U666 ( .A(n1), .ZN(n9) );
  INV_X1 U667 ( .A(n1), .ZN(n10) );
  INV_X1 U668 ( .A(n1), .ZN(n11) );
  CLKBUF_X1 U669 ( .A(n264), .Z(n12) );
  CLKBUF_X1 U670 ( .A(n264), .Z(n13) );
  INV_X1 U671 ( .A(n19), .ZN(n17) );
  INV_X1 U672 ( .A(n12), .ZN(n18) );
  INV_X1 U673 ( .A(n12), .ZN(n19) );
  INV_X1 U674 ( .A(n264), .ZN(n20) );
  INV_X1 U675 ( .A(n13), .ZN(n21) );
  INV_X1 U676 ( .A(n13), .ZN(n22) );
  CLKBUF_X1 U677 ( .A(n263), .Z(n23) );
  CLKBUF_X1 U678 ( .A(n263), .Z(n24) );
  CLKBUF_X1 U679 ( .A(n263), .Z(n25) );
  INV_X1 U680 ( .A(n23), .ZN(n30) );
  INV_X1 U681 ( .A(n24), .ZN(n31) );
  INV_X1 U682 ( .A(n25), .ZN(n32) );
endmodule


module PG_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module Gblock_0 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n2) );
endmodule


module Gblock_8 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_7 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_6 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_5 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_4 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_3 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_2 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module Gblock_1 ( Pik, Gik, Gk_1j, Gij );
  input Pik, Gik, Gk_1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk_1j), .A(Gik), .ZN(n3) );
endmodule


module PGblock_0 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_26 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_25 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_24 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_23 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_22 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_21 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_20 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_19 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_18 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_17 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_16 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_15 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_14 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_13 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_12 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_11 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_10 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_9 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_8 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_7 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_6 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_5 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_4 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
endmodule


module PGblock_3 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_2 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module PGblock_1 ( Pik, Gik, Pk_1j, Gk_1j, Pij, Gij );
  input Pik, Gik, Pk_1j, Gk_1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk_1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk_1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module carry_generator_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [32:1] A;
  input [32:1] B;
  output [7:0] Co;
  input Cin;
  wire   G_16__16_, G_16__15_, G_16__13_, G_16__9_, G_15__15_, G_14__14_,
         G_14__13_, G_13__13_, G_12__12_, G_12__11_, G_12__9_, G_11__11_,
         G_10__10_, G_10__9_, G_9__9_, G_8__8_, G_8__7_, G_8__5_, G_7__7_,
         G_6__6_, G_6__5_, G_5__5_, G_4__4_, G_4__3_, G_3__3_, G_2__2_,
         G_2__1_, G_1__1_, P_16__16_, P_16__15_, P_16__13_, P_16__9_,
         P_15__15_, P_14__14_, P_14__13_, P_13__13_, P_12__12_, P_12__11_,
         P_12__9_, P_11__11_, P_10__10_, P_10__9_, P_9__9_, P_8__8_, P_8__7_,
         P_8__5_, P_7__7_, P_6__6_, P_6__5_, P_5__5_, P_4__4_, P_4__3_,
         P_3__3_, P_2__2_, G_32__32_, G_32__31_, G_32__29_, G_32__25_,
         G_32__17_, G_31__31_, G_30__30_, G_30__29_, G_29__29_, G_28__28_,
         G_28__27_, G_28__25_, G_28__17_, G_27__27_, G_26__26_, G_26__25_,
         G_25__25_, G_24__24_, G_24__23_, G_24__21_, G_24__17_, G_23__23_,
         G_22__22_, G_22__21_, G_21__21_, G_20__20_, G_20__19_, G_20__17_,
         G_19__19_, G_18__18_, G_18__17_, G_17__17_, P_32__32_, P_32__31_,
         P_32__29_, P_32__25_, P_32__17_, P_31__31_, P_30__30_, P_30__29_,
         P_29__29_, P_28__28_, P_28__27_, P_28__25_, P_28__17_, P_27__27_,
         P_26__26_, P_26__25_, P_25__25_, P_24__24_, P_24__23_, P_24__21_,
         P_24__17_, P_23__23_, P_22__22_, P_22__21_, P_21__21_, P_20__20_,
         P_20__19_, P_20__17_, P_19__19_, P_18__18_, P_18__17_, P_17__17_, n3,
         n1, n2;

  PG_net_0 PGnetblock_2 ( .a(A[2]), .b(B[2]), .p(P_2__2_), .g(G_2__2_) );
  PG_net_30 PGnetblock_3 ( .a(A[3]), .b(B[3]), .p(P_3__3_), .g(G_3__3_) );
  PG_net_29 PGnetblock_4 ( .a(A[4]), .b(B[4]), .p(P_4__4_), .g(G_4__4_) );
  PG_net_28 PGnetblock_5 ( .a(A[5]), .b(B[5]), .p(P_5__5_), .g(G_5__5_) );
  PG_net_27 PGnetblock_6 ( .a(A[6]), .b(B[6]), .p(P_6__6_), .g(G_6__6_) );
  PG_net_26 PGnetblock_7 ( .a(A[7]), .b(B[7]), .p(P_7__7_), .g(G_7__7_) );
  PG_net_25 PGnetblock_8 ( .a(A[8]), .b(B[8]), .p(P_8__8_), .g(G_8__8_) );
  PG_net_24 PGnetblock_9 ( .a(A[9]), .b(B[9]), .p(P_9__9_), .g(G_9__9_) );
  PG_net_23 PGnetblock_10 ( .a(A[10]), .b(B[10]), .p(P_10__10_), .g(G_10__10_)
         );
  PG_net_22 PGnetblock_11 ( .a(A[11]), .b(B[11]), .p(P_11__11_), .g(G_11__11_)
         );
  PG_net_21 PGnetblock_12 ( .a(A[12]), .b(B[12]), .p(P_12__12_), .g(G_12__12_)
         );
  PG_net_20 PGnetblock_13 ( .a(A[13]), .b(B[13]), .p(P_13__13_), .g(G_13__13_)
         );
  PG_net_19 PGnetblock_14 ( .a(A[14]), .b(B[14]), .p(P_14__14_), .g(G_14__14_)
         );
  PG_net_18 PGnetblock_15 ( .a(A[15]), .b(B[15]), .p(P_15__15_), .g(G_15__15_)
         );
  PG_net_17 PGnetblock_16 ( .a(A[16]), .b(B[16]), .p(P_16__16_), .g(G_16__16_)
         );
  PG_net_16 PGnetblock_17 ( .a(A[17]), .b(B[17]), .p(P_17__17_), .g(G_17__17_)
         );
  PG_net_15 PGnetblock_18 ( .a(A[18]), .b(B[18]), .p(P_18__18_), .g(G_18__18_)
         );
  PG_net_14 PGnetblock_19 ( .a(A[19]), .b(B[19]), .p(P_19__19_), .g(G_19__19_)
         );
  PG_net_13 PGnetblock_20 ( .a(A[20]), .b(B[20]), .p(P_20__20_), .g(G_20__20_)
         );
  PG_net_12 PGnetblock_21 ( .a(A[21]), .b(B[21]), .p(P_21__21_), .g(G_21__21_)
         );
  PG_net_11 PGnetblock_22 ( .a(A[22]), .b(B[22]), .p(P_22__22_), .g(G_22__22_)
         );
  PG_net_10 PGnetblock_23 ( .a(A[23]), .b(B[23]), .p(P_23__23_), .g(G_23__23_)
         );
  PG_net_9 PGnetblock_24 ( .a(A[24]), .b(B[24]), .p(P_24__24_), .g(G_24__24_)
         );
  PG_net_8 PGnetblock_25 ( .a(A[25]), .b(B[25]), .p(P_25__25_), .g(G_25__25_)
         );
  PG_net_7 PGnetblock_26 ( .a(A[26]), .b(B[26]), .p(P_26__26_), .g(G_26__26_)
         );
  PG_net_6 PGnetblock_27 ( .a(A[27]), .b(B[27]), .p(P_27__27_), .g(G_27__27_)
         );
  PG_net_5 PGnetblock_28 ( .a(A[28]), .b(B[28]), .p(P_28__28_), .g(G_28__28_)
         );
  PG_net_4 PGnetblock_29 ( .a(A[29]), .b(B[29]), .p(P_29__29_), .g(G_29__29_)
         );
  PG_net_3 PGnetblock_30 ( .a(A[30]), .b(B[30]), .p(P_30__30_), .g(G_30__30_)
         );
  PG_net_2 PGnetblock_31 ( .a(A[31]), .b(B[31]), .p(P_31__31_), .g(G_31__31_)
         );
  PG_net_1 PGnetblock_32 ( .a(A[32]), .b(B[32]), .p(P_32__32_), .g(G_32__32_)
         );
  Gblock_0 GB_low_1_2 ( .Pik(P_2__2_), .Gik(G_2__2_), .Gk_1j(G_1__1_), .Gij(
        G_2__1_) );
  Gblock_8 GB_low_2_4 ( .Pik(P_4__3_), .Gik(G_4__3_), .Gk_1j(G_2__1_), .Gij(
        Co[0]) );
  Gblock_7 GB_low_3_8 ( .Pik(P_8__5_), .Gik(G_8__5_), .Gk_1j(Co[0]), .Gij(
        Co[1]) );
  Gblock_6 GB_high_4_16_0 ( .Pik(P_16__9_), .Gik(G_16__9_), .Gk_1j(Co[1]), 
        .Gij(Co[3]) );
  Gblock_5 GB_high_4_16_1 ( .Pik(P_12__9_), .Gik(G_12__9_), .Gk_1j(Co[1]), 
        .Gij(Co[2]) );
  Gblock_4 GB_high_5_32_0 ( .Pik(P_32__17_), .Gik(G_32__17_), .Gk_1j(Co[3]), 
        .Gij(Co[7]) );
  Gblock_3 GB_high_5_32_1 ( .Pik(P_28__17_), .Gik(G_28__17_), .Gk_1j(Co[3]), 
        .Gij(Co[6]) );
  Gblock_2 GB_high_5_32_2 ( .Pik(P_24__17_), .Gik(G_24__17_), .Gk_1j(Co[3]), 
        .Gij(Co[5]) );
  Gblock_1 GB_high_5_32_3 ( .Pik(P_20__17_), .Gik(G_20__17_), .Gk_1j(Co[3]), 
        .Gij(Co[4]) );
  PGblock_0 PGB_low_1_4 ( .Pik(P_4__4_), .Gik(G_4__4_), .Pk_1j(P_3__3_), 
        .Gk_1j(G_3__3_), .Pij(P_4__3_), .Gij(G_4__3_) );
  PGblock_26 PGB_low_1_6 ( .Pik(P_6__6_), .Gik(G_6__6_), .Pk_1j(P_5__5_), 
        .Gk_1j(G_5__5_), .Pij(P_6__5_), .Gij(G_6__5_) );
  PGblock_25 PGB_low_1_8 ( .Pik(P_8__8_), .Gik(G_8__8_), .Pk_1j(P_7__7_), 
        .Gk_1j(G_7__7_), .Pij(P_8__7_), .Gij(G_8__7_) );
  PGblock_24 PGB_low_1_10 ( .Pik(P_10__10_), .Gik(G_10__10_), .Pk_1j(P_9__9_), 
        .Gk_1j(G_9__9_), .Pij(P_10__9_), .Gij(G_10__9_) );
  PGblock_23 PGB_low_1_12 ( .Pik(P_12__12_), .Gik(G_12__12_), .Pk_1j(P_11__11_), .Gk_1j(G_11__11_), .Pij(P_12__11_), .Gij(G_12__11_) );
  PGblock_22 PGB_low_1_14 ( .Pik(P_14__14_), .Gik(G_14__14_), .Pk_1j(P_13__13_), .Gk_1j(G_13__13_), .Pij(P_14__13_), .Gij(G_14__13_) );
  PGblock_21 PGB_low_1_16 ( .Pik(P_16__16_), .Gik(G_16__16_), .Pk_1j(P_15__15_), .Gk_1j(G_15__15_), .Pij(P_16__15_), .Gij(G_16__15_) );
  PGblock_20 PGB_low_1_18 ( .Pik(P_18__18_), .Gik(G_18__18_), .Pk_1j(P_17__17_), .Gk_1j(G_17__17_), .Pij(P_18__17_), .Gij(G_18__17_) );
  PGblock_19 PGB_low_1_20 ( .Pik(P_20__20_), .Gik(G_20__20_), .Pk_1j(P_19__19_), .Gk_1j(G_19__19_), .Pij(P_20__19_), .Gij(G_20__19_) );
  PGblock_18 PGB_low_1_22 ( .Pik(P_22__22_), .Gik(G_22__22_), .Pk_1j(P_21__21_), .Gk_1j(G_21__21_), .Pij(P_22__21_), .Gij(G_22__21_) );
  PGblock_17 PGB_low_1_24 ( .Pik(P_24__24_), .Gik(G_24__24_), .Pk_1j(P_23__23_), .Gk_1j(G_23__23_), .Pij(P_24__23_), .Gij(G_24__23_) );
  PGblock_16 PGB_low_1_26 ( .Pik(P_26__26_), .Gik(G_26__26_), .Pk_1j(P_25__25_), .Gk_1j(G_25__25_), .Pij(P_26__25_), .Gij(G_26__25_) );
  PGblock_15 PGB_low_1_28 ( .Pik(P_28__28_), .Gik(G_28__28_), .Pk_1j(P_27__27_), .Gk_1j(G_27__27_), .Pij(P_28__27_), .Gij(G_28__27_) );
  PGblock_14 PGB_low_1_30 ( .Pik(P_30__30_), .Gik(G_30__30_), .Pk_1j(P_29__29_), .Gk_1j(G_29__29_), .Pij(P_30__29_), .Gij(G_30__29_) );
  PGblock_13 PGB_low_1_32 ( .Pik(P_32__32_), .Gik(G_32__32_), .Pk_1j(P_31__31_), .Gk_1j(G_31__31_), .Pij(P_32__31_), .Gij(G_32__31_) );
  PGblock_12 PGB_low_2_8 ( .Pik(P_8__7_), .Gik(G_8__7_), .Pk_1j(P_6__5_), 
        .Gk_1j(G_6__5_), .Pij(P_8__5_), .Gij(G_8__5_) );
  PGblock_11 PGB_low_2_12 ( .Pik(P_12__11_), .Gik(G_12__11_), .Pk_1j(P_10__9_), 
        .Gk_1j(G_10__9_), .Pij(P_12__9_), .Gij(G_12__9_) );
  PGblock_10 PGB_low_2_16 ( .Pik(P_16__15_), .Gik(G_16__15_), .Pk_1j(P_14__13_), .Gk_1j(G_14__13_), .Pij(P_16__13_), .Gij(G_16__13_) );
  PGblock_9 PGB_low_2_20 ( .Pik(P_20__19_), .Gik(G_20__19_), .Pk_1j(P_18__17_), 
        .Gk_1j(G_18__17_), .Pij(P_20__17_), .Gij(G_20__17_) );
  PGblock_8 PGB_low_2_24 ( .Pik(P_24__23_), .Gik(G_24__23_), .Pk_1j(P_22__21_), 
        .Gk_1j(G_22__21_), .Pij(P_24__21_), .Gij(G_24__21_) );
  PGblock_7 PGB_low_2_28 ( .Pik(P_28__27_), .Gik(G_28__27_), .Pk_1j(P_26__25_), 
        .Gk_1j(G_26__25_), .Pij(P_28__25_), .Gij(G_28__25_) );
  PGblock_6 PGB_low_2_32 ( .Pik(P_32__31_), .Gik(G_32__31_), .Pk_1j(P_30__29_), 
        .Gk_1j(G_30__29_), .Pij(P_32__29_), .Gij(G_32__29_) );
  PGblock_5 PGB_low_3_16 ( .Pik(P_16__13_), .Gik(G_16__13_), .Pk_1j(P_12__9_), 
        .Gk_1j(G_12__9_), .Pij(P_16__9_), .Gij(G_16__9_) );
  PGblock_4 PGB_low_3_24 ( .Pik(P_24__21_), .Gik(G_24__21_), .Pk_1j(P_20__17_), 
        .Gk_1j(G_20__17_), .Pij(P_24__17_), .Gij(G_24__17_) );
  PGblock_3 PGB_low_3_32 ( .Pik(P_32__29_), .Gik(G_32__29_), .Pk_1j(P_28__25_), 
        .Gk_1j(G_28__25_), .Pij(P_32__25_), .Gij(G_32__25_) );
  PGblock_2 PGB_high_4_32_0 ( .Pik(P_32__25_), .Gik(G_32__25_), .Pk_1j(
        P_24__17_), .Gk_1j(G_24__17_), .Pij(P_32__17_), .Gij(G_32__17_) );
  PGblock_1 PGB_high_4_32_1 ( .Pik(P_28__25_), .Gik(G_28__25_), .Pk_1j(
        P_24__17_), .Gk_1j(G_24__17_), .Pij(P_28__17_), .Gij(G_28__17_) );
  INV_X1 U1 ( .A(A[1]), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(G_1__1_) );
  INV_X1 U3 ( .A(B[1]), .ZN(n2) );
  OAI21_X1 U4 ( .B1(A[1]), .B2(B[1]), .A(Cin), .ZN(n3) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_0 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n6, n7, n8, n9, n5;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n6), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n6) );
  INV_X1 U6 ( .A(n8), .ZN(S[1]) );
  AOI22_X1 U7 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n8) );
  INV_X1 U8 ( .A(n7), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n7) );
  INV_X1 U10 ( .A(n9), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n9) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_7 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_6 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_5 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_4 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_3 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_2 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U5 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U7 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U8 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U9 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module carry_select_basic_N4_1 ( A, B, C_i, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_i;
  wire   n5, n10, n11, n12, n13;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  RCA_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(Y1) );
  RCA_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(Y2) );
  INV_X1 U3 ( .A(C_i), .ZN(n5) );
  INV_X1 U4 ( .A(n13), .ZN(S[3]) );
  AOI22_X1 U5 ( .A1(Y1[3]), .A2(n5), .B1(Y2[3]), .B2(C_i), .ZN(n13) );
  INV_X1 U6 ( .A(n11), .ZN(S[1]) );
  AOI22_X1 U7 ( .A1(Y1[1]), .A2(n5), .B1(Y2[1]), .B2(C_i), .ZN(n11) );
  INV_X1 U8 ( .A(n12), .ZN(S[2]) );
  AOI22_X1 U9 ( .A1(Y1[2]), .A2(n5), .B1(Y2[2]), .B2(C_i), .ZN(n12) );
  INV_X1 U10 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U11 ( .A1(Y1[0]), .A2(n5), .B1(Y2[0]), .B2(C_i), .ZN(n10) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  carry_select_basic_N4_0 CSBI_1 ( .A(A[3:0]), .B(B[3:0]), .C_i(Ci[0]), .S(
        S[3:0]) );
  carry_select_basic_N4_7 CSBI_2 ( .A(A[7:4]), .B(B[7:4]), .C_i(Ci[1]), .S(
        S[7:4]) );
  carry_select_basic_N4_6 CSBI_3 ( .A(A[11:8]), .B(B[11:8]), .C_i(Ci[2]), .S(
        S[11:8]) );
  carry_select_basic_N4_5 CSBI_4 ( .A(A[15:12]), .B(B[15:12]), .C_i(Ci[3]), 
        .S(S[15:12]) );
  carry_select_basic_N4_4 CSBI_5 ( .A(A[19:16]), .B(B[19:16]), .C_i(Ci[4]), 
        .S(S[19:16]) );
  carry_select_basic_N4_3 CSBI_6 ( .A(A[23:20]), .B(B[23:20]), .C_i(Ci[5]), 
        .S(S[23:20]) );
  carry_select_basic_N4_2 CSBI_7 ( .A(A[27:24]), .B(B[27:24]), .C_i(Ci[6]), 
        .S(S[27:24]) );
  carry_select_basic_N4_1 CSBI_8 ( .A(A[31:28]), .B(B[31:28]), .C_i(Ci[7]), 
        .S(S[31:28]) );
endmodule


module P4Adder_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [7:1] Csum;

  carry_generator_NBIT32_NBIT_PER_BLOCK4 Carrygen0 ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Csum}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 Sumgen0 ( .A(A), .B(B), .Ci({Csum, 
        Cin}), .S(S) );
endmodule


module booth_encoder_numBit16 ( B, SEL_out );
  input [15:0] B;
  output [23:0] SEL_out;

  assign SEL_out[0] = 1'b0;
  assign SEL_out[23] = B[15];
  assign SEL_out[22] = B[14];
  assign SEL_out[20] = B[13];
  assign SEL_out[21] = B[13];
  assign SEL_out[19] = B[12];
  assign SEL_out[17] = B[11];
  assign SEL_out[18] = B[11];
  assign SEL_out[16] = B[10];
  assign SEL_out[14] = B[9];
  assign SEL_out[15] = B[9];
  assign SEL_out[13] = B[8];
  assign SEL_out[11] = B[7];
  assign SEL_out[12] = B[7];
  assign SEL_out[10] = B[6];
  assign SEL_out[8] = B[5];
  assign SEL_out[9] = B[5];
  assign SEL_out[7] = B[4];
  assign SEL_out[5] = B[3];
  assign SEL_out[6] = B[3];
  assign SEL_out[4] = B[2];
  assign SEL_out[2] = B[1];
  assign SEL_out[3] = B[1];
  assign SEL_out[1] = B[0];

endmodule


module mux5to1_numBit32_0 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  OAI33_X1 U109 ( .A1(n91), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n90), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n8) );
  BUF_X1 U2 ( .A(n10), .Z(n4) );
  BUF_X1 U3 ( .A(n10), .Z(n77) );
  BUF_X1 U4 ( .A(n10), .Z(n78) );
  INV_X1 U5 ( .A(SEL_in[1]), .ZN(n90) );
  AOI222_X1 U6 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n68) );
  AOI222_X1 U7 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n66) );
  AOI222_X1 U8 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n64) );
  AOI222_X1 U9 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n62) );
  AOI222_X1 U10 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n60) );
  AOI222_X1 U11 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n58) );
  AOI222_X1 U12 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n56) );
  AOI222_X1 U13 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n54) );
  AOI222_X1 U14 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n52) );
  AOI222_X1 U15 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n50) );
  AOI222_X1 U16 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n48) );
  AOI222_X1 U17 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n46) );
  AOI222_X1 U18 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n44) );
  AOI222_X1 U19 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n42) );
  AOI222_X1 U20 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n22) );
  AOI222_X1 U21 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n20) );
  AOI222_X1 U22 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n18) );
  AOI222_X1 U23 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n16) );
  AOI222_X1 U24 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n14) );
  AOI222_X1 U25 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n12) );
  AOI222_X1 U26 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n70) );
  AOI222_X1 U27 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n40) );
  AOI222_X1 U28 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n38) );
  AOI222_X1 U29 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n36) );
  AOI222_X1 U30 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n34) );
  AOI222_X1 U31 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n32) );
  AOI222_X1 U32 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n30) );
  AOI222_X1 U33 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n28) );
  AOI222_X1 U34 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n26) );
  AOI222_X1 U35 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n24) );
  BUF_X1 U36 ( .A(n9), .Z(n79) );
  BUF_X1 U37 ( .A(n9), .Z(n80) );
  BUF_X1 U38 ( .A(n7), .Z(n85) );
  BUF_X1 U39 ( .A(n7), .Z(n86) );
  BUF_X1 U40 ( .A(n89), .Z(n1) );
  BUF_X1 U41 ( .A(n89), .Z(n2) );
  NOR2_X1 U42 ( .A1(n88), .A2(n75), .ZN(n10) );
  INV_X1 U43 ( .A(n74), .ZN(n88) );
  BUF_X1 U44 ( .A(n89), .Z(n3) );
  BUF_X1 U45 ( .A(n9), .Z(n81) );
  BUF_X1 U46 ( .A(n7), .Z(n87) );
  NOR4_X1 U47 ( .A1(n76), .A2(n85), .A3(n79), .A4(n82), .ZN(n74) );
  NOR3_X1 U48 ( .A1(n90), .A2(SEL_in[2]), .A3(n91), .ZN(n7) );
  BUF_X1 U49 ( .A(n8), .Z(n82) );
  BUF_X1 U50 ( .A(n8), .Z(n83) );
  BUF_X1 U51 ( .A(n8), .Z(n84) );
  NOR2_X1 U52 ( .A1(n90), .A2(n91), .ZN(n75) );
  AND3_X1 U53 ( .A1(n91), .A2(n90), .A3(SEL_in[2]), .ZN(n9) );
  NAND2_X1 U54 ( .A1(n65), .A2(n66), .ZN(Z[3]) );
  INV_X1 U55 ( .A(n73), .ZN(n89) );
  AOI21_X1 U56 ( .B1(n74), .B2(n75), .A(n76), .ZN(n73) );
  AOI22_X1 U57 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n69) );
  AOI22_X1 U58 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n67) );
  AOI22_X1 U59 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n65) );
  AOI22_X1 U60 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n63) );
  AOI22_X1 U61 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n61) );
  AOI22_X1 U62 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n59) );
  AOI22_X1 U63 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n57) );
  AOI22_X1 U64 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n55) );
  AOI22_X1 U65 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n53) );
  AOI22_X1 U66 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n51) );
  AOI22_X1 U67 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n49) );
  AOI22_X1 U68 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n47) );
  AOI22_X1 U69 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n45) );
  AOI22_X1 U70 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n43) );
  NOR3_X1 U71 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n76) );
  AOI222_X1 U72 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n72) );
  AOI22_X1 U73 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n41) );
  AOI22_X1 U74 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n23) );
  AOI22_X1 U75 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n21) );
  AOI22_X1 U76 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n19) );
  AOI22_X1 U77 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n17) );
  AOI22_X1 U78 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n15) );
  AOI22_X1 U79 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n13) );
  AOI22_X1 U80 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n11) );
  AOI22_X1 U81 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n71) );
  AOI22_X1 U82 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n33) );
  AOI22_X1 U83 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n31) );
  AOI22_X1 U84 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n29) );
  AOI22_X1 U85 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n27) );
  AOI22_X1 U86 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n25) );
  NAND2_X1 U87 ( .A1(n63), .A2(n64), .ZN(Z[4]) );
  NAND2_X1 U88 ( .A1(n61), .A2(n62), .ZN(Z[5]) );
  NAND2_X1 U89 ( .A1(n59), .A2(n60), .ZN(Z[6]) );
  NAND2_X1 U90 ( .A1(n57), .A2(n58), .ZN(Z[7]) );
  NAND2_X1 U91 ( .A1(n55), .A2(n56), .ZN(Z[8]) );
  NAND2_X1 U92 ( .A1(n53), .A2(n54), .ZN(Z[9]) );
  NAND2_X1 U93 ( .A1(n51), .A2(n52), .ZN(Z[10]) );
  NAND2_X1 U94 ( .A1(n49), .A2(n50), .ZN(Z[11]) );
  NAND2_X1 U95 ( .A1(n47), .A2(n48), .ZN(Z[12]) );
  NAND2_X1 U96 ( .A1(n45), .A2(n46), .ZN(Z[13]) );
  NAND2_X1 U97 ( .A1(n43), .A2(n44), .ZN(Z[14]) );
  NAND2_X1 U98 ( .A1(n41), .A2(n42), .ZN(Z[15]) );
  NAND2_X1 U99 ( .A1(n39), .A2(n40), .ZN(Z[16]) );
  AOI22_X1 U100 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n39) );
  NAND2_X1 U101 ( .A1(n37), .A2(n38), .ZN(Z[17]) );
  AOI22_X1 U102 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n37) );
  NAND2_X1 U103 ( .A1(n35), .A2(n36), .ZN(Z[18]) );
  AOI22_X1 U104 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n35) );
  NAND2_X1 U105 ( .A1(n33), .A2(n34), .ZN(Z[19]) );
  NAND2_X1 U106 ( .A1(n31), .A2(n32), .ZN(Z[20]) );
  NAND2_X1 U107 ( .A1(n29), .A2(n30), .ZN(Z[21]) );
  NAND2_X1 U108 ( .A1(n27), .A2(n28), .ZN(Z[22]) );
  NAND2_X1 U110 ( .A1(n25), .A2(n26), .ZN(Z[23]) );
  NAND2_X1 U111 ( .A1(n23), .A2(n24), .ZN(Z[24]) );
  NAND2_X1 U112 ( .A1(n21), .A2(n22), .ZN(Z[25]) );
  NAND2_X1 U113 ( .A1(n19), .A2(n20), .ZN(Z[26]) );
  NAND2_X1 U114 ( .A1(n17), .A2(n18), .ZN(Z[27]) );
  NAND2_X1 U115 ( .A1(n15), .A2(n16), .ZN(Z[28]) );
  NAND2_X1 U116 ( .A1(n13), .A2(n14), .ZN(Z[29]) );
  NAND2_X1 U117 ( .A1(n11), .A2(n12), .ZN(Z[30]) );
  NAND2_X1 U118 ( .A1(n67), .A2(n68), .ZN(Z[2]) );
  NAND2_X1 U119 ( .A1(n71), .A2(n72), .ZN(Z[0]) );
  NAND2_X1 U120 ( .A1(n69), .A2(n70), .ZN(Z[1]) );
  NAND2_X1 U121 ( .A1(n5), .A2(n6), .ZN(Z[31]) );
  AOI22_X1 U122 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n5) );
  AOI222_X1 U123 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n6) );
  INV_X1 U124 ( .A(SEL_in[0]), .ZN(n91) );
endmodule


module mux5to1_numBit32_7 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  AOI222_X1 U6 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  AOI222_X1 U7 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  AOI222_X1 U8 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  AOI222_X1 U9 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  AOI222_X1 U10 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  AOI222_X1 U11 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  AOI222_X1 U12 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  AOI222_X1 U13 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  AOI222_X1 U14 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  AOI222_X1 U15 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  AOI222_X1 U16 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  AOI222_X1 U17 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  BUF_X1 U18 ( .A(n89), .Z(n1) );
  BUF_X1 U19 ( .A(n89), .Z(n2) );
  NOR2_X1 U20 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U21 ( .A(n94), .ZN(n88) );
  BUF_X1 U22 ( .A(n89), .Z(n3) );
  NOR4_X1 U23 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U24 ( .A(n160), .Z(n82) );
  BUF_X1 U25 ( .A(n160), .Z(n83) );
  BUF_X1 U26 ( .A(n159), .Z(n79) );
  BUF_X1 U27 ( .A(n159), .Z(n80) );
  BUF_X1 U28 ( .A(n161), .Z(n85) );
  BUF_X1 U29 ( .A(n161), .Z(n86) );
  BUF_X1 U30 ( .A(n160), .Z(n84) );
  NOR2_X1 U31 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U32 ( .A(n159), .Z(n81) );
  BUF_X1 U33 ( .A(n161), .Z(n87) );
  INV_X1 U34 ( .A(n95), .ZN(n89) );
  AOI21_X1 U35 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  AOI222_X1 U36 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  AOI222_X1 U37 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  AOI222_X1 U38 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  AOI222_X1 U39 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  AOI222_X1 U40 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  AOI222_X1 U41 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  AOI222_X1 U42 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  AOI222_X1 U43 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  AOI222_X1 U44 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  AOI222_X1 U45 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  AOI222_X1 U46 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  AOI222_X1 U47 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  AOI222_X1 U48 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  AOI222_X1 U49 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NOR3_X1 U50 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U51 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U52 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U53 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U54 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U55 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI222_X1 U56 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  AOI22_X1 U57 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI22_X1 U58 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U59 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  AOI22_X1 U60 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI22_X1 U61 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  NAND2_X1 U62 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U63 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  NAND2_X1 U64 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U65 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  NAND2_X1 U66 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U67 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  NAND2_X1 U68 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U69 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  NAND2_X1 U70 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U71 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  NAND2_X1 U72 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U73 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  NAND2_X1 U74 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U75 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  NAND2_X1 U76 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U77 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  NAND2_X1 U78 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U79 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  NAND2_X1 U80 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U81 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  NAND2_X1 U82 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U83 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  NAND2_X1 U84 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U85 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  NAND2_X1 U86 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  NAND2_X1 U87 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  NAND2_X1 U88 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  NAND2_X1 U89 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U90 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  NAND2_X1 U91 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U92 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  NAND2_X1 U93 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U94 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  NAND2_X1 U95 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U96 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  NAND2_X1 U97 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U98 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  NAND2_X1 U99 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U100 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  NAND2_X1 U101 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U102 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  NAND2_X1 U103 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U104 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  NAND2_X1 U105 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U106 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  NAND2_X1 U107 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U108 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  NAND2_X1 U110 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U111 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  NAND2_X1 U112 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U113 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  NAND2_X1 U114 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U115 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  NAND2_X1 U116 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U117 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  NAND2_X1 U118 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U119 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  NAND2_X1 U120 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U121 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U122 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
  AOI222_X1 U123 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  AOI222_X1 U124 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
endmodule


module mux5to1_numBit32_6 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI222_X1 U30 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  AOI22_X1 U31 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  NAND2_X1 U32 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U33 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U34 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U35 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U36 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U37 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U38 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U39 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U40 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U41 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U42 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U43 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U44 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U45 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U46 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U47 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U48 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U49 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U50 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U51 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U52 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U53 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U54 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U55 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U56 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U57 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U58 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U59 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U60 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U61 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U62 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U63 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U64 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U65 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U66 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U67 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U68 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U69 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U70 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U71 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U72 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U73 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U74 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U75 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U76 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U77 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U78 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U79 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U80 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U81 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U82 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U83 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U84 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U85 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U86 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U87 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U88 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U89 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U90 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U91 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U92 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U93 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U94 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U95 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U96 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U97 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U98 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U99 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U100 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), .C2(n81), .ZN(n152) );
  NAND2_X1 U101 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U102 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U103 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), .C2(n81), .ZN(n154) );
  NAND2_X1 U104 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U105 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U106 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), .C2(n81), .ZN(n156) );
  NAND2_X1 U107 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U108 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U110 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U111 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U112 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U113 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U114 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U115 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U116 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U117 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U118 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U119 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U120 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U121 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U122 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_5 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U26 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI222_X1 U29 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  AOI22_X1 U30 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  NAND2_X1 U31 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U33 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U35 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U36 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U37 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U38 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U39 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U40 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U41 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U42 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U43 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U44 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U45 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U46 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U47 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U48 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U49 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U50 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U51 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U52 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U53 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U54 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U55 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U56 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U57 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U58 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U59 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U60 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U61 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U62 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U63 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U64 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U65 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U66 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U67 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U68 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U69 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U70 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U71 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U72 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U73 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U74 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U75 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U76 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U77 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U78 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U79 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U80 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U81 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U82 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U83 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U84 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U85 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U86 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U87 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U88 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U89 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U90 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U91 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U92 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U93 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U94 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U95 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U96 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U97 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U98 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U99 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U100 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U101 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U102 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U103 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U104 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U105 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U106 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U107 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U108 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U110 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U111 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U112 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U113 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U114 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U115 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U116 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U117 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U118 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U119 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U120 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U121 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module mux5to1_numBit32_4 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI222_X1 U30 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  AOI22_X1 U31 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  NAND2_X1 U32 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U33 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U34 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U35 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U36 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U37 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  NAND2_X1 U38 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U39 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U40 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U41 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U43 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U44 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U45 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U46 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U47 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U48 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U49 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U50 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U51 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U52 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U53 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U54 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U55 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U56 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U57 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U58 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U59 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U60 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U61 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U62 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U63 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U64 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U65 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U66 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U67 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U68 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U69 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U70 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U71 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U72 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U73 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U74 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U75 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U76 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U77 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U78 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U79 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U80 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U81 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U82 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U83 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U84 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U85 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U86 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U87 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U88 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U89 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U90 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U91 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U92 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U93 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U94 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U95 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U96 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U97 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U98 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U99 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U100 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U101 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U102 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U103 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U104 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U105 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U106 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U107 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U108 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U110 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U111 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U112 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U113 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U114 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U115 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U116 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U117 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U118 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U119 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U120 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U121 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U122 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_3 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n91), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n90), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n90), .A2(n91), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n90), .A2(SEL_in[2]), .A3(n91), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n91) );
  AND3_X1 U26 ( .A1(n91), .A2(n90), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n90) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI222_X1 U29 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), 
        .C2(n79), .ZN(n118) );
  AOI22_X1 U30 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  NAND2_X1 U31 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U32 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U33 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U34 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U35 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U36 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  NAND2_X1 U37 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U38 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U39 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U40 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U41 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U42 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U43 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U44 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U45 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U46 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U47 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U48 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U49 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U50 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U51 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U52 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U53 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U54 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U55 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U57 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U58 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U59 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U60 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U61 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U62 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U63 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U64 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U65 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U66 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U67 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U68 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U69 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U70 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U71 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U72 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U73 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U74 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U75 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U76 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U77 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U78 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U79 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U80 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U81 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U82 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U83 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U84 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U85 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U86 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U87 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U88 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U89 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U90 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), 
        .C2(n79), .ZN(n116) );
  NAND2_X1 U91 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U92 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U93 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U94 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U95 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U96 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U97 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U98 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U99 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U100 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U101 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U102 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U103 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U104 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U105 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U106 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U107 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U108 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U110 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U111 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U112 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U113 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U114 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U115 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U116 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U117 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U118 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U119 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U120 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U121 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module mux5to1_numBit32_2 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  AOI222_X1 U5 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), 
        .C2(n81), .ZN(n162) );
  BUF_X1 U6 ( .A(n89), .Z(n1) );
  BUF_X1 U7 ( .A(n89), .Z(n2) );
  NOR2_X1 U8 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U9 ( .A(n94), .ZN(n88) );
  BUF_X1 U10 ( .A(n89), .Z(n3) );
  NOR4_X1 U11 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U12 ( .A(n160), .Z(n82) );
  BUF_X1 U13 ( .A(n160), .Z(n83) );
  BUF_X1 U14 ( .A(n159), .Z(n79) );
  BUF_X1 U15 ( .A(n159), .Z(n80) );
  BUF_X1 U16 ( .A(n161), .Z(n85) );
  BUF_X1 U17 ( .A(n161), .Z(n86) );
  BUF_X1 U18 ( .A(n160), .Z(n84) );
  NOR2_X1 U19 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U20 ( .A(n159), .Z(n81) );
  BUF_X1 U21 ( .A(n161), .Z(n87) );
  INV_X1 U22 ( .A(n95), .ZN(n89) );
  AOI21_X1 U23 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U24 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U25 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U26 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U27 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U28 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U29 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI222_X1 U30 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), 
        .C2(n80), .ZN(n122) );
  AOI22_X1 U31 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  NAND2_X1 U32 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U33 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U34 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U35 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI22_X1 U36 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  AOI222_X1 U37 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  NAND2_X1 U38 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U39 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U40 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U41 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U42 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U43 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U44 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U45 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U46 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U47 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U48 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U49 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U50 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U51 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U52 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U53 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U54 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U55 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U56 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U57 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U58 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U59 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U60 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U61 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U62 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U63 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U64 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U65 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U67 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U68 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U69 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U70 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U71 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U72 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U73 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U74 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U75 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U76 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U77 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U78 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U79 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U80 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U81 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U82 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U83 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U84 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U85 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), 
        .C2(n80), .ZN(n120) );
  NAND2_X1 U86 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U87 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U88 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U89 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U90 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U91 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U92 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U93 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U94 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U95 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U96 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U97 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U98 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U99 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U100 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U101 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U102 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U103 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U104 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U105 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U106 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U107 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U108 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U110 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U111 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U112 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U113 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U114 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U115 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U116 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U117 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U118 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U119 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), .C2(n79), .ZN(n116) );
  NAND2_X1 U120 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U121 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U122 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), .C2(n79), .ZN(n118) );
  NAND2_X1 U123 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U124 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
endmodule


module mux5to1_numBit32_1 ( IN1, IN2, IN3, IN4, IN5, SEL_in, Z );
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [2:0] SEL_in;
  output [31:0] Z;
  wire   n1, n2, n3, n4, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  OAI33_X1 U109 ( .A1(n90), .A2(SEL_in[2]), .A3(SEL_in[1]), .B1(n91), .B2(
        SEL_in[2]), .B3(SEL_in[0]), .ZN(n160) );
  BUF_X1 U2 ( .A(n158), .Z(n4) );
  BUF_X1 U3 ( .A(n158), .Z(n77) );
  BUF_X1 U4 ( .A(n158), .Z(n78) );
  BUF_X1 U5 ( .A(n89), .Z(n1) );
  BUF_X1 U6 ( .A(n89), .Z(n2) );
  NOR2_X1 U7 ( .A1(n88), .A2(n93), .ZN(n158) );
  INV_X1 U8 ( .A(n94), .ZN(n88) );
  BUF_X1 U9 ( .A(n89), .Z(n3) );
  NOR4_X1 U10 ( .A1(n92), .A2(n85), .A3(n79), .A4(n82), .ZN(n94) );
  BUF_X1 U11 ( .A(n160), .Z(n82) );
  BUF_X1 U12 ( .A(n160), .Z(n83) );
  BUF_X1 U13 ( .A(n159), .Z(n79) );
  BUF_X1 U14 ( .A(n159), .Z(n80) );
  BUF_X1 U15 ( .A(n161), .Z(n85) );
  BUF_X1 U16 ( .A(n161), .Z(n86) );
  BUF_X1 U17 ( .A(n160), .Z(n84) );
  NOR2_X1 U18 ( .A1(n91), .A2(n90), .ZN(n93) );
  BUF_X1 U19 ( .A(n159), .Z(n81) );
  BUF_X1 U20 ( .A(n161), .Z(n87) );
  INV_X1 U21 ( .A(n95), .ZN(n89) );
  AOI21_X1 U22 ( .B1(n94), .B2(n93), .A(n92), .ZN(n95) );
  NOR3_X1 U23 ( .A1(n91), .A2(SEL_in[2]), .A3(n90), .ZN(n161) );
  NOR3_X1 U24 ( .A1(SEL_in[1]), .A2(SEL_in[2]), .A3(SEL_in[0]), .ZN(n92) );
  INV_X1 U25 ( .A(SEL_in[0]), .ZN(n90) );
  AND3_X1 U26 ( .A1(n90), .A2(n91), .A3(SEL_in[2]), .ZN(n159) );
  INV_X1 U27 ( .A(SEL_in[1]), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n127), .A2(n126), .ZN(Z[15]) );
  AOI222_X1 U29 ( .A1(IN4[15]), .A2(n86), .B1(IN2[15]), .B2(n83), .C1(IN5[15]), 
        .C2(n80), .ZN(n126) );
  AOI22_X1 U30 ( .A1(IN3[15]), .A2(n77), .B1(IN1[15]), .B2(n2), .ZN(n127) );
  NAND2_X1 U31 ( .A1(n129), .A2(n128), .ZN(Z[16]) );
  AOI22_X1 U32 ( .A1(IN3[16]), .A2(n77), .B1(IN1[16]), .B2(n2), .ZN(n129) );
  AOI222_X1 U33 ( .A1(IN4[16]), .A2(n86), .B1(IN2[16]), .B2(n83), .C1(IN5[16]), 
        .C2(n80), .ZN(n128) );
  NAND2_X1 U34 ( .A1(n131), .A2(n130), .ZN(Z[17]) );
  AOI22_X1 U35 ( .A1(IN3[17]), .A2(n77), .B1(IN1[17]), .B2(n2), .ZN(n131) );
  AOI222_X1 U36 ( .A1(IN4[17]), .A2(n86), .B1(IN2[17]), .B2(n83), .C1(IN5[17]), 
        .C2(n80), .ZN(n130) );
  NAND2_X1 U37 ( .A1(n133), .A2(n132), .ZN(Z[18]) );
  AOI22_X1 U38 ( .A1(IN3[18]), .A2(n77), .B1(IN1[18]), .B2(n2), .ZN(n133) );
  AOI222_X1 U39 ( .A1(IN4[18]), .A2(n86), .B1(IN2[18]), .B2(n83), .C1(IN5[18]), 
        .C2(n80), .ZN(n132) );
  NAND2_X1 U40 ( .A1(n135), .A2(n134), .ZN(Z[19]) );
  AOI22_X1 U41 ( .A1(IN3[19]), .A2(n77), .B1(IN1[19]), .B2(n2), .ZN(n135) );
  AOI222_X1 U42 ( .A1(IN4[19]), .A2(n86), .B1(IN2[19]), .B2(n83), .C1(IN5[19]), 
        .C2(n80), .ZN(n134) );
  NAND2_X1 U43 ( .A1(n137), .A2(n136), .ZN(Z[20]) );
  AOI22_X1 U44 ( .A1(IN3[20]), .A2(n77), .B1(IN1[20]), .B2(n2), .ZN(n137) );
  AOI222_X1 U45 ( .A1(IN4[20]), .A2(n86), .B1(IN2[20]), .B2(n83), .C1(IN5[20]), 
        .C2(n80), .ZN(n136) );
  NAND2_X1 U46 ( .A1(n139), .A2(n138), .ZN(Z[21]) );
  AOI22_X1 U47 ( .A1(IN3[21]), .A2(n77), .B1(IN1[21]), .B2(n2), .ZN(n139) );
  AOI222_X1 U48 ( .A1(IN4[21]), .A2(n86), .B1(IN2[21]), .B2(n83), .C1(IN5[21]), 
        .C2(n80), .ZN(n138) );
  NAND2_X1 U49 ( .A1(n141), .A2(n140), .ZN(Z[22]) );
  AOI22_X1 U50 ( .A1(IN3[22]), .A2(n77), .B1(IN1[22]), .B2(n2), .ZN(n141) );
  AOI222_X1 U51 ( .A1(IN4[22]), .A2(n86), .B1(IN2[22]), .B2(n83), .C1(IN5[22]), 
        .C2(n80), .ZN(n140) );
  NAND2_X1 U52 ( .A1(n143), .A2(n142), .ZN(Z[23]) );
  AOI22_X1 U53 ( .A1(IN3[23]), .A2(n77), .B1(IN1[23]), .B2(n2), .ZN(n143) );
  AOI222_X1 U54 ( .A1(IN4[23]), .A2(n86), .B1(IN2[23]), .B2(n83), .C1(IN5[23]), 
        .C2(n80), .ZN(n142) );
  NAND2_X1 U55 ( .A1(n145), .A2(n144), .ZN(Z[24]) );
  AOI22_X1 U56 ( .A1(IN3[24]), .A2(n78), .B1(IN1[24]), .B2(n3), .ZN(n145) );
  AOI222_X1 U57 ( .A1(IN4[24]), .A2(n86), .B1(IN2[24]), .B2(n83), .C1(IN5[24]), 
        .C2(n80), .ZN(n144) );
  NAND2_X1 U58 ( .A1(n147), .A2(n146), .ZN(Z[25]) );
  AOI22_X1 U59 ( .A1(IN3[25]), .A2(n78), .B1(IN1[25]), .B2(n3), .ZN(n147) );
  AOI222_X1 U60 ( .A1(IN4[25]), .A2(n87), .B1(IN2[25]), .B2(n84), .C1(IN5[25]), 
        .C2(n81), .ZN(n146) );
  NAND2_X1 U61 ( .A1(n149), .A2(n148), .ZN(Z[26]) );
  AOI22_X1 U62 ( .A1(IN3[26]), .A2(n78), .B1(IN1[26]), .B2(n3), .ZN(n149) );
  AOI222_X1 U63 ( .A1(IN4[26]), .A2(n87), .B1(IN2[26]), .B2(n84), .C1(IN5[26]), 
        .C2(n81), .ZN(n148) );
  NAND2_X1 U64 ( .A1(n151), .A2(n150), .ZN(Z[27]) );
  AOI22_X1 U65 ( .A1(IN3[27]), .A2(n78), .B1(IN1[27]), .B2(n3), .ZN(n151) );
  AOI222_X1 U66 ( .A1(IN4[27]), .A2(n87), .B1(IN2[27]), .B2(n84), .C1(IN5[27]), 
        .C2(n81), .ZN(n150) );
  NAND2_X1 U67 ( .A1(n153), .A2(n152), .ZN(Z[28]) );
  AOI22_X1 U68 ( .A1(IN3[28]), .A2(n78), .B1(IN1[28]), .B2(n3), .ZN(n153) );
  AOI222_X1 U69 ( .A1(IN4[28]), .A2(n87), .B1(IN2[28]), .B2(n84), .C1(IN5[28]), 
        .C2(n81), .ZN(n152) );
  NAND2_X1 U70 ( .A1(n155), .A2(n154), .ZN(Z[29]) );
  AOI22_X1 U71 ( .A1(IN3[29]), .A2(n78), .B1(IN1[29]), .B2(n3), .ZN(n155) );
  AOI222_X1 U72 ( .A1(IN4[29]), .A2(n87), .B1(IN2[29]), .B2(n84), .C1(IN5[29]), 
        .C2(n81), .ZN(n154) );
  NAND2_X1 U73 ( .A1(n157), .A2(n156), .ZN(Z[30]) );
  AOI22_X1 U74 ( .A1(IN3[30]), .A2(n78), .B1(IN1[30]), .B2(n3), .ZN(n157) );
  AOI222_X1 U75 ( .A1(IN4[30]), .A2(n87), .B1(IN2[30]), .B2(n84), .C1(IN5[30]), 
        .C2(n81), .ZN(n156) );
  NAND2_X1 U76 ( .A1(n125), .A2(n124), .ZN(Z[14]) );
  AOI22_X1 U77 ( .A1(IN3[14]), .A2(n77), .B1(IN1[14]), .B2(n2), .ZN(n125) );
  AOI222_X1 U78 ( .A1(IN4[14]), .A2(n86), .B1(IN2[14]), .B2(n83), .C1(IN5[14]), 
        .C2(n80), .ZN(n124) );
  NAND2_X1 U79 ( .A1(n97), .A2(n96), .ZN(Z[0]) );
  AOI22_X1 U80 ( .A1(IN3[0]), .A2(n4), .B1(IN1[0]), .B2(n1), .ZN(n97) );
  AOI222_X1 U81 ( .A1(IN4[0]), .A2(n85), .B1(IN2[0]), .B2(n82), .C1(IN5[0]), 
        .C2(n79), .ZN(n96) );
  NAND2_X1 U82 ( .A1(n99), .A2(n98), .ZN(Z[1]) );
  AOI22_X1 U83 ( .A1(IN3[1]), .A2(n4), .B1(IN1[1]), .B2(n1), .ZN(n99) );
  AOI222_X1 U84 ( .A1(IN4[1]), .A2(n85), .B1(IN2[1]), .B2(n82), .C1(IN5[1]), 
        .C2(n79), .ZN(n98) );
  NAND2_X1 U85 ( .A1(n101), .A2(n100), .ZN(Z[2]) );
  AOI22_X1 U86 ( .A1(IN3[2]), .A2(n4), .B1(IN1[2]), .B2(n1), .ZN(n101) );
  AOI222_X1 U87 ( .A1(IN4[2]), .A2(n85), .B1(IN2[2]), .B2(n82), .C1(IN5[2]), 
        .C2(n79), .ZN(n100) );
  NAND2_X1 U88 ( .A1(n103), .A2(n102), .ZN(Z[3]) );
  AOI22_X1 U89 ( .A1(IN3[3]), .A2(n4), .B1(IN1[3]), .B2(n1), .ZN(n103) );
  AOI222_X1 U90 ( .A1(IN4[3]), .A2(n85), .B1(IN2[3]), .B2(n82), .C1(IN5[3]), 
        .C2(n79), .ZN(n102) );
  NAND2_X1 U91 ( .A1(n105), .A2(n104), .ZN(Z[4]) );
  AOI22_X1 U92 ( .A1(IN3[4]), .A2(n4), .B1(IN1[4]), .B2(n1), .ZN(n105) );
  AOI222_X1 U93 ( .A1(IN4[4]), .A2(n85), .B1(IN2[4]), .B2(n82), .C1(IN5[4]), 
        .C2(n79), .ZN(n104) );
  NAND2_X1 U94 ( .A1(n107), .A2(n106), .ZN(Z[5]) );
  AOI22_X1 U95 ( .A1(IN3[5]), .A2(n4), .B1(IN1[5]), .B2(n1), .ZN(n107) );
  AOI222_X1 U96 ( .A1(IN4[5]), .A2(n85), .B1(IN2[5]), .B2(n82), .C1(IN5[5]), 
        .C2(n79), .ZN(n106) );
  NAND2_X1 U97 ( .A1(n109), .A2(n108), .ZN(Z[6]) );
  AOI22_X1 U98 ( .A1(IN3[6]), .A2(n4), .B1(IN1[6]), .B2(n1), .ZN(n109) );
  AOI222_X1 U99 ( .A1(IN4[6]), .A2(n85), .B1(IN2[6]), .B2(n82), .C1(IN5[6]), 
        .C2(n79), .ZN(n108) );
  NAND2_X1 U100 ( .A1(n111), .A2(n110), .ZN(Z[7]) );
  AOI22_X1 U101 ( .A1(IN3[7]), .A2(n4), .B1(IN1[7]), .B2(n1), .ZN(n111) );
  AOI222_X1 U102 ( .A1(IN4[7]), .A2(n85), .B1(IN2[7]), .B2(n82), .C1(IN5[7]), 
        .C2(n79), .ZN(n110) );
  NAND2_X1 U103 ( .A1(n113), .A2(n112), .ZN(Z[8]) );
  AOI22_X1 U104 ( .A1(IN3[8]), .A2(n4), .B1(IN1[8]), .B2(n1), .ZN(n113) );
  AOI222_X1 U105 ( .A1(IN4[8]), .A2(n85), .B1(IN2[8]), .B2(n82), .C1(IN5[8]), 
        .C2(n79), .ZN(n112) );
  NAND2_X1 U106 ( .A1(n115), .A2(n114), .ZN(Z[9]) );
  AOI22_X1 U107 ( .A1(IN3[9]), .A2(n4), .B1(IN1[9]), .B2(n1), .ZN(n115) );
  AOI222_X1 U108 ( .A1(IN4[9]), .A2(n85), .B1(IN2[9]), .B2(n82), .C1(IN5[9]), 
        .C2(n79), .ZN(n114) );
  NAND2_X1 U110 ( .A1(n117), .A2(n116), .ZN(Z[10]) );
  AOI22_X1 U111 ( .A1(IN3[10]), .A2(n4), .B1(IN1[10]), .B2(n1), .ZN(n117) );
  AOI222_X1 U112 ( .A1(IN4[10]), .A2(n85), .B1(IN2[10]), .B2(n82), .C1(IN5[10]), .C2(n79), .ZN(n116) );
  NAND2_X1 U113 ( .A1(n119), .A2(n118), .ZN(Z[11]) );
  AOI22_X1 U114 ( .A1(IN3[11]), .A2(n4), .B1(IN1[11]), .B2(n1), .ZN(n119) );
  AOI222_X1 U115 ( .A1(IN4[11]), .A2(n85), .B1(IN2[11]), .B2(n82), .C1(IN5[11]), .C2(n79), .ZN(n118) );
  NAND2_X1 U116 ( .A1(n121), .A2(n120), .ZN(Z[12]) );
  AOI22_X1 U117 ( .A1(IN3[12]), .A2(n77), .B1(IN1[12]), .B2(n2), .ZN(n121) );
  AOI222_X1 U118 ( .A1(IN4[12]), .A2(n86), .B1(IN2[12]), .B2(n83), .C1(IN5[12]), .C2(n80), .ZN(n120) );
  NAND2_X1 U119 ( .A1(n123), .A2(n122), .ZN(Z[13]) );
  AOI22_X1 U120 ( .A1(IN3[13]), .A2(n77), .B1(IN1[13]), .B2(n2), .ZN(n123) );
  AOI222_X1 U121 ( .A1(IN4[13]), .A2(n86), .B1(IN2[13]), .B2(n83), .C1(IN5[13]), .C2(n80), .ZN(n122) );
  NAND2_X1 U122 ( .A1(n163), .A2(n162), .ZN(Z[31]) );
  AOI22_X1 U123 ( .A1(IN3[31]), .A2(n78), .B1(IN1[31]), .B2(n3), .ZN(n163) );
  AOI222_X1 U124 ( .A1(IN4[31]), .A2(n87), .B1(IN2[31]), .B2(n84), .C1(IN5[31]), .C2(n81), .ZN(n162) );
endmodule


module rca_bhv_numBit32_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_0 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_0_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_6 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_6_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_5 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_5_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_4 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_4_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_3 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_3_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_2 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_2_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module rca_bhv_numBit32_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module rca_bhv_numBit32_1 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;


  rca_bhv_numBit32_1_DW01_add_0 add_1_root_add_35_2 ( .A({A[31], A}), .B({
        B[31], B}), .CI(Ci), .SUM({Co, S}) );
endmodule


module BOOTHMUL_numBit16 ( A, B, P );
  input [15:0] A;
  input [15:0] B;
  output [31:0] P;
  wire   rca_out_5__31_, rca_out_5__30_, rca_out_5__29_, rca_out_5__28_,
         rca_out_5__27_, rca_out_5__26_, rca_out_5__25_, rca_out_5__24_,
         rca_out_5__23_, rca_out_5__22_, rca_out_5__21_, rca_out_5__20_,
         rca_out_5__19_, rca_out_5__18_, rca_out_5__17_, rca_out_5__16_,
         rca_out_5__15_, rca_out_5__14_, rca_out_5__13_, rca_out_5__12_,
         rca_out_5__11_, rca_out_5__10_, rca_out_5__9_, rca_out_5__8_,
         rca_out_5__7_, rca_out_5__6_, rca_out_5__5_, rca_out_5__4_,
         rca_out_5__3_, rca_out_5__2_, rca_out_5__1_, rca_out_5__0_,
         rca_out_4__31_, rca_out_4__30_, rca_out_4__29_, rca_out_4__28_,
         rca_out_4__27_, rca_out_4__26_, rca_out_4__25_, rca_out_4__24_,
         rca_out_4__23_, rca_out_4__22_, rca_out_4__21_, rca_out_4__20_,
         rca_out_4__19_, rca_out_4__18_, rca_out_4__17_, rca_out_4__16_,
         rca_out_4__15_, rca_out_4__14_, rca_out_4__13_, rca_out_4__12_,
         rca_out_4__11_, rca_out_4__10_, rca_out_4__9_, rca_out_4__8_,
         rca_out_4__7_, rca_out_4__6_, rca_out_4__5_, rca_out_4__4_,
         rca_out_4__3_, rca_out_4__2_, rca_out_4__1_, rca_out_4__0_,
         rca_out_3__31_, rca_out_3__30_, rca_out_3__29_, rca_out_3__28_,
         rca_out_3__27_, rca_out_3__26_, rca_out_3__25_, rca_out_3__24_,
         rca_out_3__23_, rca_out_3__22_, rca_out_3__21_, rca_out_3__20_,
         rca_out_3__19_, rca_out_3__18_, rca_out_3__17_, rca_out_3__16_,
         rca_out_3__15_, rca_out_3__14_, rca_out_3__13_, rca_out_3__12_,
         rca_out_3__11_, rca_out_3__10_, rca_out_3__9_, rca_out_3__8_,
         rca_out_3__7_, rca_out_3__6_, rca_out_3__5_, rca_out_3__4_,
         rca_out_3__3_, rca_out_3__2_, rca_out_3__1_, rca_out_3__0_,
         rca_out_2__31_, rca_out_2__30_, rca_out_2__29_, rca_out_2__28_,
         rca_out_2__27_, rca_out_2__26_, rca_out_2__25_, rca_out_2__24_,
         rca_out_2__23_, rca_out_2__22_, rca_out_2__21_, rca_out_2__20_,
         rca_out_2__19_, rca_out_2__18_, rca_out_2__17_, rca_out_2__16_,
         rca_out_2__15_, rca_out_2__14_, rca_out_2__13_, rca_out_2__12_,
         rca_out_2__11_, rca_out_2__10_, rca_out_2__9_, rca_out_2__8_,
         rca_out_2__7_, rca_out_2__6_, rca_out_2__5_, rca_out_2__4_,
         rca_out_2__3_, rca_out_2__2_, rca_out_2__1_, rca_out_2__0_,
         rca_out_1__31_, rca_out_1__30_, rca_out_1__29_, rca_out_1__28_,
         rca_out_1__27_, rca_out_1__26_, rca_out_1__25_, rca_out_1__24_,
         rca_out_1__23_, rca_out_1__22_, rca_out_1__21_, rca_out_1__20_,
         rca_out_1__19_, rca_out_1__18_, rca_out_1__17_, rca_out_1__16_,
         rca_out_1__15_, rca_out_1__14_, rca_out_1__13_, rca_out_1__12_,
         rca_out_1__11_, rca_out_1__10_, rca_out_1__9_, rca_out_1__8_,
         rca_out_1__7_, rca_out_1__6_, rca_out_1__5_, rca_out_1__4_,
         rca_out_1__3_, rca_out_1__2_, rca_out_1__1_, rca_out_1__0_,
         rca_out_0__31_, rca_out_0__30_, rca_out_0__29_, rca_out_0__28_,
         rca_out_0__27_, rca_out_0__26_, rca_out_0__25_, rca_out_0__24_,
         rca_out_0__23_, rca_out_0__22_, rca_out_0__21_, rca_out_0__20_,
         rca_out_0__19_, rca_out_0__18_, rca_out_0__17_, rca_out_0__16_,
         rca_out_0__15_, rca_out_0__14_, rca_out_0__13_, rca_out_0__12_,
         rca_out_0__11_, rca_out_0__10_, rca_out_0__9_, rca_out_0__8_,
         rca_out_0__7_, rca_out_0__6_, rca_out_0__5_, rca_out_0__4_,
         rca_out_0__3_, rca_out_0__2_, rca_out_0__1_, rca_out_0__0_,
         add_65_carry_2_, add_65_carry_3_, add_65_carry_4_, add_65_carry_5_,
         add_65_carry_6_, add_65_carry_7_, add_65_carry_8_, add_65_carry_9_,
         add_65_carry_10_, add_65_carry_11_, add_65_carry_12_,
         add_65_carry_13_, add_65_carry_14_, add_65_carry_15_, add_65_A_0_,
         add_65_A_1_, add_65_A_2_, add_65_A_3_, add_65_A_4_, add_65_A_5_,
         add_65_A_6_, add_65_A_7_, add_65_A_8_, add_65_A_9_, add_65_A_10_,
         add_65_A_11_, add_65_A_12_, add_65_A_13_, add_65_A_14_, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, SYNOPSYS_UNCONNECTED_1;
  wire   [23:0] encoder_out;
  wire   [31:0] A_minus;
  wire   [255:0] sum_op;

  booth_encoder_numBit16 encode ( .B(B), .SEL_out({encoder_out[23:1], 
        SYNOPSYS_UNCONNECTED_1}) );
  mux5to1_numBit32_0 mux0_0 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n48, n48, n49, n48, n48, n49, n48, n49, n48, n48, n48, 
        n49, n48, n49, n48, n49, n48, A[14:0]}), .IN3({n35, n31, n31, n36, n31, 
        n35, n31, n36, n31, n36, n32, n35, n32, n35, n33, n34, A_minus[15], n2, 
        n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, 
        A_minus[0]}), .IN4({n42, n42, n42, n42, n42, n42, n42, n42, n42, n42, 
        n42, n43, n43, n43, n43, n43, A[14:0], 1'b0}), .IN5({n41, n41, n41, 
        n41, n41, n41, n40, n40, n39, n40, n38, n39, n38, n38, n39, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0}), .SEL_in({encoder_out[2:1], 1'b0}), .Z(
        sum_op[31:0]) );
  mux5to1_numBit32_7 mux_i_1 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n51, n51, n51, n51, n51, n50, n50, n50, n50, n50, 
        n49, n49, n49, n49, A[14:0], 1'b0, 1'b0}), .IN3({n31, n36, n31, n35, 
        n31, n35, n32, n36, n32, n35, n33, n34, n33, n34, A_minus[15], n2, n4, 
        n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 
        1'b0, 1'b0}), .IN4({n47, n47, n47, n47, n46, n47, n47, n47, n46, n46, 
        n46, n46, n46, n42, A[14:0], 1'b0, 1'b0, 1'b0}), .IN5({n41, n41, n40, 
        n40, n40, n40, n40, n41, n37, n39, n37, n39, n37, A_minus[15], n2, n4, 
        n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 
        1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[5:3]), .Z(sum_op[63:32]) );
  mux5to1_numBit32_6 mux_i_2 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({A[15], A[15], A[15], A[15], A[15], A[15], n48, A[15], 
        A[15], n53, n53, n53, n53, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({
        n31, n36, n31, n36, n32, n36, n32, n36, n33, n34, n33, n34, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n46, n46, n46, 
        n46, n46, n47, n46, n47, n45, n47, n47, n47, A[14:0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN5({n41, n41, n40, n40, n39, n39, n38, n38, n37, n37, 
        n38, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, 
        n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[8:6]), .Z(sum_op[95:64]) );
  mux5to1_numBit32_5 mux_i_3 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n52, n50, n53, n53, n53, n53, n53, n53, n53, n53, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n31, n35, n32, 
        n35, n32, n36, n33, n34, n33, n34, A_minus[15], n2, n4, n6, n8, n10, 
        n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n45, n45, n45, n45, n45, n45, n45, n45, 
        n45, n45, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({
        n40, n40, n39, n39, n37, n38, n38, n37, n38, A_minus[15], n2, n4, n6, 
        n8, n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[11:9]), .Z(
        sum_op[127:96]) );
  mux5to1_numBit32_4 mux_i_4 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n52, n52, n52, n52, n52, n52, n52, n52, n52, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n31, n36, n32, 
        n36, n33, n34, n33, n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, 
        n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n44, n44, n44, n44, n44, n44, n44, n44, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5(
        {n39, n39, n38, n41, n37, n38, n39, A_minus[15], n2, n4, n6, n8, n10, 
        n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(encoder_out[14:12]), .Z(sum_op[159:128]) );
  mux5to1_numBit32_3 mux_i_5 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n51, n51, n51, n51, n51, n51, n51, A[14:0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n32, n35, n32, 
        n35, n33, n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, 
        n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n43, n44, n44, n44, n44, 
        A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN5({n40, n39, n37, n38, n37, A_minus[15], n2, n4, n6, n8, 
        n10, n12, n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[17:15]), .Z(sum_op[191:160]) );
  mux5to1_numBit32_2 mux_i_6 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n50, n50, n50, n50, n50, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n32, n35, n33, 
        n34, A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, 
        n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n43, n43, n43, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN5({n37, n38, n37, A_minus[15], n2, n4, n6, n8, n10, n12, 
        n14, n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL_in(
        encoder_out[20:18]), .Z(sum_op[223:192]) );
  mux5to1_numBit32_1 mux_i_7 ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN2({n49, n49, n50, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({n33, n34, 
        A_minus[15], n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, 
        n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({n43, n45, A[14:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN5({n37, A_minus[15], n2, n4, n6, n8, n10, n12, n14, 
        n16, n18, n20, n22, n24, n26, n28, A_minus[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL_in(encoder_out[23:21]), .Z(sum_op[255:224]) );
  rca_bhv_numBit32_0 rca0_0 ( .A(sum_op[31:0]), .B(sum_op[63:32]), .Ci(1'b0), 
        .S({rca_out_0__31_, rca_out_0__30_, rca_out_0__29_, rca_out_0__28_, 
        rca_out_0__27_, rca_out_0__26_, rca_out_0__25_, rca_out_0__24_, 
        rca_out_0__23_, rca_out_0__22_, rca_out_0__21_, rca_out_0__20_, 
        rca_out_0__19_, rca_out_0__18_, rca_out_0__17_, rca_out_0__16_, 
        rca_out_0__15_, rca_out_0__14_, rca_out_0__13_, rca_out_0__12_, 
        rca_out_0__11_, rca_out_0__10_, rca_out_0__9_, rca_out_0__8_, 
        rca_out_0__7_, rca_out_0__6_, rca_out_0__5_, rca_out_0__4_, 
        rca_out_0__3_, rca_out_0__2_, rca_out_0__1_, rca_out_0__0_}) );
  rca_bhv_numBit32_6 rca_i_1 ( .A({rca_out_0__31_, rca_out_0__30_, 
        rca_out_0__29_, rca_out_0__28_, rca_out_0__27_, rca_out_0__26_, 
        rca_out_0__25_, rca_out_0__24_, rca_out_0__23_, rca_out_0__22_, 
        rca_out_0__21_, rca_out_0__20_, rca_out_0__19_, rca_out_0__18_, 
        rca_out_0__17_, rca_out_0__16_, rca_out_0__15_, rca_out_0__14_, 
        rca_out_0__13_, rca_out_0__12_, rca_out_0__11_, rca_out_0__10_, 
        rca_out_0__9_, rca_out_0__8_, rca_out_0__7_, rca_out_0__6_, 
        rca_out_0__5_, rca_out_0__4_, rca_out_0__3_, rca_out_0__2_, 
        rca_out_0__1_, rca_out_0__0_}), .B(sum_op[95:64]), .Ci(1'b0), .S({
        rca_out_1__31_, rca_out_1__30_, rca_out_1__29_, rca_out_1__28_, 
        rca_out_1__27_, rca_out_1__26_, rca_out_1__25_, rca_out_1__24_, 
        rca_out_1__23_, rca_out_1__22_, rca_out_1__21_, rca_out_1__20_, 
        rca_out_1__19_, rca_out_1__18_, rca_out_1__17_, rca_out_1__16_, 
        rca_out_1__15_, rca_out_1__14_, rca_out_1__13_, rca_out_1__12_, 
        rca_out_1__11_, rca_out_1__10_, rca_out_1__9_, rca_out_1__8_, 
        rca_out_1__7_, rca_out_1__6_, rca_out_1__5_, rca_out_1__4_, 
        rca_out_1__3_, rca_out_1__2_, rca_out_1__1_, rca_out_1__0_}) );
  rca_bhv_numBit32_5 rca_i_2 ( .A({rca_out_1__31_, rca_out_1__30_, 
        rca_out_1__29_, rca_out_1__28_, rca_out_1__27_, rca_out_1__26_, 
        rca_out_1__25_, rca_out_1__24_, rca_out_1__23_, rca_out_1__22_, 
        rca_out_1__21_, rca_out_1__20_, rca_out_1__19_, rca_out_1__18_, 
        rca_out_1__17_, rca_out_1__16_, rca_out_1__15_, rca_out_1__14_, 
        rca_out_1__13_, rca_out_1__12_, rca_out_1__11_, rca_out_1__10_, 
        rca_out_1__9_, rca_out_1__8_, rca_out_1__7_, rca_out_1__6_, 
        rca_out_1__5_, rca_out_1__4_, rca_out_1__3_, rca_out_1__2_, 
        rca_out_1__1_, rca_out_1__0_}), .B(sum_op[127:96]), .Ci(1'b0), .S({
        rca_out_2__31_, rca_out_2__30_, rca_out_2__29_, rca_out_2__28_, 
        rca_out_2__27_, rca_out_2__26_, rca_out_2__25_, rca_out_2__24_, 
        rca_out_2__23_, rca_out_2__22_, rca_out_2__21_, rca_out_2__20_, 
        rca_out_2__19_, rca_out_2__18_, rca_out_2__17_, rca_out_2__16_, 
        rca_out_2__15_, rca_out_2__14_, rca_out_2__13_, rca_out_2__12_, 
        rca_out_2__11_, rca_out_2__10_, rca_out_2__9_, rca_out_2__8_, 
        rca_out_2__7_, rca_out_2__6_, rca_out_2__5_, rca_out_2__4_, 
        rca_out_2__3_, rca_out_2__2_, rca_out_2__1_, rca_out_2__0_}) );
  rca_bhv_numBit32_4 rca_i_3 ( .A({rca_out_2__31_, rca_out_2__30_, 
        rca_out_2__29_, rca_out_2__28_, rca_out_2__27_, rca_out_2__26_, 
        rca_out_2__25_, rca_out_2__24_, rca_out_2__23_, rca_out_2__22_, 
        rca_out_2__21_, rca_out_2__20_, rca_out_2__19_, rca_out_2__18_, 
        rca_out_2__17_, rca_out_2__16_, rca_out_2__15_, rca_out_2__14_, 
        rca_out_2__13_, rca_out_2__12_, rca_out_2__11_, rca_out_2__10_, 
        rca_out_2__9_, rca_out_2__8_, rca_out_2__7_, rca_out_2__6_, 
        rca_out_2__5_, rca_out_2__4_, rca_out_2__3_, rca_out_2__2_, 
        rca_out_2__1_, rca_out_2__0_}), .B(sum_op[159:128]), .Ci(1'b0), .S({
        rca_out_3__31_, rca_out_3__30_, rca_out_3__29_, rca_out_3__28_, 
        rca_out_3__27_, rca_out_3__26_, rca_out_3__25_, rca_out_3__24_, 
        rca_out_3__23_, rca_out_3__22_, rca_out_3__21_, rca_out_3__20_, 
        rca_out_3__19_, rca_out_3__18_, rca_out_3__17_, rca_out_3__16_, 
        rca_out_3__15_, rca_out_3__14_, rca_out_3__13_, rca_out_3__12_, 
        rca_out_3__11_, rca_out_3__10_, rca_out_3__9_, rca_out_3__8_, 
        rca_out_3__7_, rca_out_3__6_, rca_out_3__5_, rca_out_3__4_, 
        rca_out_3__3_, rca_out_3__2_, rca_out_3__1_, rca_out_3__0_}) );
  rca_bhv_numBit32_3 rca_i_4 ( .A({rca_out_3__31_, rca_out_3__30_, 
        rca_out_3__29_, rca_out_3__28_, rca_out_3__27_, rca_out_3__26_, 
        rca_out_3__25_, rca_out_3__24_, rca_out_3__23_, rca_out_3__22_, 
        rca_out_3__21_, rca_out_3__20_, rca_out_3__19_, rca_out_3__18_, 
        rca_out_3__17_, rca_out_3__16_, rca_out_3__15_, rca_out_3__14_, 
        rca_out_3__13_, rca_out_3__12_, rca_out_3__11_, rca_out_3__10_, 
        rca_out_3__9_, rca_out_3__8_, rca_out_3__7_, rca_out_3__6_, 
        rca_out_3__5_, rca_out_3__4_, rca_out_3__3_, rca_out_3__2_, 
        rca_out_3__1_, rca_out_3__0_}), .B(sum_op[191:160]), .Ci(1'b0), .S({
        rca_out_4__31_, rca_out_4__30_, rca_out_4__29_, rca_out_4__28_, 
        rca_out_4__27_, rca_out_4__26_, rca_out_4__25_, rca_out_4__24_, 
        rca_out_4__23_, rca_out_4__22_, rca_out_4__21_, rca_out_4__20_, 
        rca_out_4__19_, rca_out_4__18_, rca_out_4__17_, rca_out_4__16_, 
        rca_out_4__15_, rca_out_4__14_, rca_out_4__13_, rca_out_4__12_, 
        rca_out_4__11_, rca_out_4__10_, rca_out_4__9_, rca_out_4__8_, 
        rca_out_4__7_, rca_out_4__6_, rca_out_4__5_, rca_out_4__4_, 
        rca_out_4__3_, rca_out_4__2_, rca_out_4__1_, rca_out_4__0_}) );
  rca_bhv_numBit32_2 rca_i_5 ( .A({rca_out_4__31_, rca_out_4__30_, 
        rca_out_4__29_, rca_out_4__28_, rca_out_4__27_, rca_out_4__26_, 
        rca_out_4__25_, rca_out_4__24_, rca_out_4__23_, rca_out_4__22_, 
        rca_out_4__21_, rca_out_4__20_, rca_out_4__19_, rca_out_4__18_, 
        rca_out_4__17_, rca_out_4__16_, rca_out_4__15_, rca_out_4__14_, 
        rca_out_4__13_, rca_out_4__12_, rca_out_4__11_, rca_out_4__10_, 
        rca_out_4__9_, rca_out_4__8_, rca_out_4__7_, rca_out_4__6_, 
        rca_out_4__5_, rca_out_4__4_, rca_out_4__3_, rca_out_4__2_, 
        rca_out_4__1_, rca_out_4__0_}), .B(sum_op[223:192]), .Ci(1'b0), .S({
        rca_out_5__31_, rca_out_5__30_, rca_out_5__29_, rca_out_5__28_, 
        rca_out_5__27_, rca_out_5__26_, rca_out_5__25_, rca_out_5__24_, 
        rca_out_5__23_, rca_out_5__22_, rca_out_5__21_, rca_out_5__20_, 
        rca_out_5__19_, rca_out_5__18_, rca_out_5__17_, rca_out_5__16_, 
        rca_out_5__15_, rca_out_5__14_, rca_out_5__13_, rca_out_5__12_, 
        rca_out_5__11_, rca_out_5__10_, rca_out_5__9_, rca_out_5__8_, 
        rca_out_5__7_, rca_out_5__6_, rca_out_5__5_, rca_out_5__4_, 
        rca_out_5__3_, rca_out_5__2_, rca_out_5__1_, rca_out_5__0_}) );
  rca_bhv_numBit32_1 rca_i_6 ( .A({rca_out_5__31_, rca_out_5__30_, 
        rca_out_5__29_, rca_out_5__28_, rca_out_5__27_, rca_out_5__26_, 
        rca_out_5__25_, rca_out_5__24_, rca_out_5__23_, rca_out_5__22_, 
        rca_out_5__21_, rca_out_5__20_, rca_out_5__19_, rca_out_5__18_, 
        rca_out_5__17_, rca_out_5__16_, rca_out_5__15_, rca_out_5__14_, 
        rca_out_5__13_, rca_out_5__12_, rca_out_5__11_, rca_out_5__10_, 
        rca_out_5__9_, rca_out_5__8_, rca_out_5__7_, rca_out_5__6_, 
        rca_out_5__5_, rca_out_5__4_, rca_out_5__3_, rca_out_5__2_, 
        rca_out_5__1_, rca_out_5__0_}), .B(sum_op[255:224]), .Ci(1'b0), .S(P)
         );
  HA_X1 add_65_U1_1_1 ( .A(add_65_A_1_), .B(add_65_A_0_), .CO(add_65_carry_2_), 
        .S(A_minus[1]) );
  HA_X1 add_65_U1_1_2 ( .A(add_65_A_2_), .B(add_65_carry_2_), .CO(
        add_65_carry_3_), .S(A_minus[2]) );
  HA_X1 add_65_U1_1_3 ( .A(add_65_A_3_), .B(add_65_carry_3_), .CO(
        add_65_carry_4_), .S(A_minus[3]) );
  HA_X1 add_65_U1_1_4 ( .A(add_65_A_4_), .B(add_65_carry_4_), .CO(
        add_65_carry_5_), .S(A_minus[4]) );
  HA_X1 add_65_U1_1_5 ( .A(add_65_A_5_), .B(add_65_carry_5_), .CO(
        add_65_carry_6_), .S(A_minus[5]) );
  HA_X1 add_65_U1_1_6 ( .A(add_65_A_6_), .B(add_65_carry_6_), .CO(
        add_65_carry_7_), .S(A_minus[6]) );
  HA_X1 add_65_U1_1_7 ( .A(add_65_A_7_), .B(add_65_carry_7_), .CO(
        add_65_carry_8_), .S(A_minus[7]) );
  HA_X1 add_65_U1_1_8 ( .A(add_65_A_8_), .B(add_65_carry_8_), .CO(
        add_65_carry_9_), .S(A_minus[8]) );
  HA_X1 add_65_U1_1_9 ( .A(add_65_A_9_), .B(add_65_carry_9_), .CO(
        add_65_carry_10_), .S(A_minus[9]) );
  HA_X1 add_65_U1_1_10 ( .A(add_65_A_10_), .B(add_65_carry_10_), .CO(
        add_65_carry_11_), .S(A_minus[10]) );
  HA_X1 add_65_U1_1_11 ( .A(add_65_A_11_), .B(add_65_carry_11_), .CO(
        add_65_carry_12_), .S(A_minus[11]) );
  HA_X1 add_65_U1_1_12 ( .A(add_65_A_12_), .B(add_65_carry_12_), .CO(
        add_65_carry_13_), .S(A_minus[12]) );
  HA_X1 add_65_U1_1_13 ( .A(add_65_A_13_), .B(add_65_carry_13_), .CO(
        add_65_carry_14_), .S(A_minus[13]) );
  HA_X1 add_65_U1_1_14 ( .A(add_65_A_14_), .B(add_65_carry_14_), .CO(
        add_65_carry_15_), .S(A_minus[14]) );
  INV_X1 U3 ( .A(A_minus[14]), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(n2) );
  INV_X1 U5 ( .A(A_minus[13]), .ZN(n3) );
  INV_X1 U6 ( .A(n3), .ZN(n4) );
  INV_X1 U7 ( .A(A_minus[12]), .ZN(n5) );
  INV_X1 U8 ( .A(n5), .ZN(n6) );
  INV_X1 U9 ( .A(A_minus[11]), .ZN(n7) );
  INV_X1 U10 ( .A(n7), .ZN(n8) );
  INV_X1 U11 ( .A(A_minus[10]), .ZN(n9) );
  INV_X1 U12 ( .A(n9), .ZN(n10) );
  INV_X1 U13 ( .A(A_minus[9]), .ZN(n11) );
  INV_X1 U14 ( .A(n11), .ZN(n12) );
  INV_X1 U15 ( .A(A_minus[8]), .ZN(n13) );
  INV_X1 U16 ( .A(n13), .ZN(n14) );
  INV_X1 U17 ( .A(A_minus[7]), .ZN(n15) );
  INV_X1 U18 ( .A(n15), .ZN(n16) );
  INV_X1 U19 ( .A(A_minus[6]), .ZN(n17) );
  INV_X1 U20 ( .A(n17), .ZN(n18) );
  INV_X1 U21 ( .A(A_minus[5]), .ZN(n19) );
  INV_X1 U22 ( .A(n19), .ZN(n20) );
  INV_X1 U23 ( .A(A_minus[4]), .ZN(n21) );
  INV_X1 U24 ( .A(n21), .ZN(n22) );
  INV_X1 U25 ( .A(A_minus[3]), .ZN(n23) );
  INV_X1 U26 ( .A(n23), .ZN(n24) );
  INV_X1 U27 ( .A(A_minus[2]), .ZN(n25) );
  INV_X1 U28 ( .A(n25), .ZN(n26) );
  INV_X1 U29 ( .A(A_minus[1]), .ZN(n27) );
  INV_X1 U30 ( .A(n27), .ZN(n28) );
  BUF_X1 U31 ( .A(n30), .Z(n40) );
  BUF_X1 U32 ( .A(n30), .Z(n39) );
  BUF_X1 U33 ( .A(n30), .Z(n37) );
  BUF_X1 U34 ( .A(n30), .Z(n38) );
  BUF_X1 U35 ( .A(n29), .Z(n36) );
  BUF_X1 U36 ( .A(n29), .Z(n31) );
  BUF_X1 U37 ( .A(n29), .Z(n33) );
  BUF_X1 U38 ( .A(n29), .Z(n35) );
  BUF_X1 U39 ( .A(n29), .Z(n32) );
  BUF_X1 U40 ( .A(n29), .Z(n34) );
  BUF_X1 U41 ( .A(n30), .Z(n41) );
  BUF_X1 U42 ( .A(A_minus[31]), .Z(n29) );
  BUF_X1 U43 ( .A(A_minus[31]), .Z(n30) );
  INV_X1 U44 ( .A(n54), .ZN(n42) );
  INV_X1 U45 ( .A(n54), .ZN(n43) );
  INV_X1 U46 ( .A(n54), .ZN(n47) );
  INV_X1 U47 ( .A(n54), .ZN(n46) );
  INV_X1 U48 ( .A(n54), .ZN(n44) );
  INV_X1 U49 ( .A(n54), .ZN(n45) );
  INV_X1 U50 ( .A(n54), .ZN(n48) );
  INV_X1 U51 ( .A(n54), .ZN(n53) );
  INV_X1 U52 ( .A(n54), .ZN(n52) );
  INV_X1 U53 ( .A(n54), .ZN(n51) );
  INV_X1 U54 ( .A(n54), .ZN(n50) );
  INV_X1 U55 ( .A(n54), .ZN(n49) );
  INV_X1 U56 ( .A(add_65_A_0_), .ZN(A_minus[0]) );
  INV_X1 U57 ( .A(A[0]), .ZN(add_65_A_0_) );
  INV_X1 U58 ( .A(A[14]), .ZN(add_65_A_14_) );
  INV_X1 U59 ( .A(A[1]), .ZN(add_65_A_1_) );
  INV_X1 U60 ( .A(A[2]), .ZN(add_65_A_2_) );
  INV_X1 U61 ( .A(A[3]), .ZN(add_65_A_3_) );
  INV_X1 U62 ( .A(A[4]), .ZN(add_65_A_4_) );
  INV_X1 U63 ( .A(A[5]), .ZN(add_65_A_5_) );
  INV_X1 U64 ( .A(A[6]), .ZN(add_65_A_6_) );
  INV_X1 U65 ( .A(A[7]), .ZN(add_65_A_7_) );
  INV_X1 U66 ( .A(A[8]), .ZN(add_65_A_8_) );
  INV_X1 U67 ( .A(A[9]), .ZN(add_65_A_9_) );
  INV_X1 U68 ( .A(A[10]), .ZN(add_65_A_10_) );
  INV_X1 U69 ( .A(A[11]), .ZN(add_65_A_11_) );
  INV_X1 U70 ( .A(A[12]), .ZN(add_65_A_12_) );
  INV_X1 U71 ( .A(A[13]), .ZN(add_65_A_13_) );
  XOR2_X2 U72 ( .A(add_65_carry_15_), .B(n54), .Z(A_minus[15]) );
  INV_X1 U73 ( .A(A[15]), .ZN(n54) );
  NOR2_X1 U74 ( .A1(add_65_carry_15_), .A2(A[15]), .ZN(A_minus[31]) );
endmodule


module mux41_NBIT32_1 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149;

  BUF_X1 U1 ( .A(n145), .Z(n72) );
  BUF_X1 U2 ( .A(n145), .Z(n73) );
  BUF_X1 U3 ( .A(n146), .Z(n75) );
  BUF_X1 U4 ( .A(n146), .Z(n76) );
  BUF_X1 U5 ( .A(n145), .Z(n74) );
  BUF_X1 U6 ( .A(n146), .Z(n77) );
  NOR2_X1 U7 ( .A1(n81), .A2(S[1]), .ZN(n145) );
  BUF_X1 U8 ( .A(n147), .Z(n78) );
  BUF_X1 U9 ( .A(n147), .Z(n79) );
  BUF_X1 U10 ( .A(n144), .Z(n1) );
  BUF_X1 U11 ( .A(n144), .Z(n70) );
  BUF_X1 U12 ( .A(n147), .Z(n80) );
  BUF_X1 U13 ( .A(n144), .Z(n71) );
  AND2_X1 U14 ( .A1(S[1]), .A2(n81), .ZN(n146) );
  NOR2_X1 U15 ( .A1(S[0]), .A2(S[1]), .ZN(n144) );
  AOI22_X1 U16 ( .A1(D[0]), .A2(n78), .B1(C[0]), .B2(n75), .ZN(n82) );
  AOI22_X1 U17 ( .A1(B[5]), .A2(n74), .B1(A[5]), .B2(n71), .ZN(n137) );
  AOI22_X1 U18 ( .A1(B[6]), .A2(n74), .B1(A[6]), .B2(n71), .ZN(n139) );
  AOI22_X1 U19 ( .A1(B[7]), .A2(n74), .B1(A[7]), .B2(n71), .ZN(n141) );
  AOI22_X1 U20 ( .A1(B[9]), .A2(n74), .B1(A[9]), .B2(n71), .ZN(n149) );
  AOI22_X1 U21 ( .A1(B[31]), .A2(n74), .B1(A[31]), .B2(n71), .ZN(n131) );
  AOI22_X1 U22 ( .A1(B[10]), .A2(n72), .B1(A[10]), .B2(n1), .ZN(n85) );
  AOI22_X1 U23 ( .A1(B[11]), .A2(n72), .B1(A[11]), .B2(n1), .ZN(n87) );
  AOI22_X1 U24 ( .A1(B[13]), .A2(n72), .B1(A[13]), .B2(n1), .ZN(n91) );
  AOI22_X1 U25 ( .A1(B[14]), .A2(n72), .B1(A[14]), .B2(n1), .ZN(n93) );
  AOI22_X1 U26 ( .A1(B[15]), .A2(n72), .B1(A[15]), .B2(n1), .ZN(n95) );
  AOI22_X1 U27 ( .A1(B[17]), .A2(n72), .B1(A[17]), .B2(n1), .ZN(n99) );
  AOI22_X1 U28 ( .A1(B[18]), .A2(n72), .B1(A[18]), .B2(n1), .ZN(n101) );
  AOI22_X1 U29 ( .A1(B[19]), .A2(n72), .B1(A[19]), .B2(n1), .ZN(n103) );
  AOI22_X1 U30 ( .A1(B[21]), .A2(n73), .B1(A[21]), .B2(n70), .ZN(n109) );
  AOI22_X1 U31 ( .A1(B[22]), .A2(n73), .B1(A[22]), .B2(n70), .ZN(n111) );
  AOI22_X1 U32 ( .A1(B[23]), .A2(n73), .B1(A[23]), .B2(n70), .ZN(n113) );
  AOI22_X1 U33 ( .A1(B[25]), .A2(n73), .B1(A[25]), .B2(n70), .ZN(n117) );
  AOI22_X1 U34 ( .A1(B[26]), .A2(n73), .B1(A[26]), .B2(n70), .ZN(n119) );
  AOI22_X1 U35 ( .A1(B[27]), .A2(n73), .B1(A[27]), .B2(n70), .ZN(n121) );
  AOI22_X1 U36 ( .A1(B[29]), .A2(n73), .B1(A[29]), .B2(n70), .ZN(n125) );
  AOI22_X1 U37 ( .A1(B[30]), .A2(n73), .B1(A[30]), .B2(n70), .ZN(n129) );
  AND2_X1 U38 ( .A1(S[1]), .A2(S[0]), .ZN(n147) );
  INV_X1 U39 ( .A(S[0]), .ZN(n81) );
  AOI22_X1 U40 ( .A1(B[3]), .A2(n74), .B1(A[3]), .B2(n71), .ZN(n133) );
  AOI22_X1 U41 ( .A1(B[4]), .A2(n74), .B1(A[4]), .B2(n71), .ZN(n135) );
  AOI22_X1 U42 ( .A1(B[8]), .A2(n74), .B1(A[8]), .B2(n71), .ZN(n143) );
  AOI22_X1 U43 ( .A1(B[1]), .A2(n72), .B1(A[1]), .B2(n1), .ZN(n105) );
  AOI22_X1 U44 ( .A1(B[2]), .A2(n73), .B1(A[2]), .B2(n70), .ZN(n127) );
  AOI22_X1 U45 ( .A1(B[12]), .A2(n72), .B1(A[12]), .B2(n1), .ZN(n89) );
  AOI22_X1 U46 ( .A1(B[16]), .A2(n72), .B1(A[16]), .B2(n1), .ZN(n97) );
  AOI22_X1 U47 ( .A1(B[20]), .A2(n73), .B1(A[20]), .B2(n70), .ZN(n107) );
  AOI22_X1 U48 ( .A1(B[24]), .A2(n73), .B1(A[24]), .B2(n70), .ZN(n115) );
  AOI22_X1 U49 ( .A1(B[28]), .A2(n73), .B1(A[28]), .B2(n70), .ZN(n123) );
  NAND2_X1 U50 ( .A1(n131), .A2(n130), .ZN(Z[31]) );
  NAND2_X1 U51 ( .A1(n83), .A2(n82), .ZN(Z[0]) );
  AOI22_X1 U52 ( .A1(B[0]), .A2(n72), .B1(A[0]), .B2(n1), .ZN(n83) );
  AOI22_X1 U53 ( .A1(D[31]), .A2(n80), .B1(C[31]), .B2(n77), .ZN(n130) );
  NAND2_X1 U54 ( .A1(n133), .A2(n132), .ZN(Z[3]) );
  AOI22_X1 U55 ( .A1(D[3]), .A2(n80), .B1(C[3]), .B2(n77), .ZN(n132) );
  NAND2_X1 U56 ( .A1(n135), .A2(n134), .ZN(Z[4]) );
  AOI22_X1 U57 ( .A1(D[4]), .A2(n80), .B1(C[4]), .B2(n77), .ZN(n134) );
  NAND2_X1 U58 ( .A1(n137), .A2(n136), .ZN(Z[5]) );
  AOI22_X1 U59 ( .A1(D[5]), .A2(n80), .B1(C[5]), .B2(n77), .ZN(n136) );
  NAND2_X1 U60 ( .A1(n139), .A2(n138), .ZN(Z[6]) );
  AOI22_X1 U61 ( .A1(D[6]), .A2(n80), .B1(C[6]), .B2(n77), .ZN(n138) );
  NAND2_X1 U62 ( .A1(n141), .A2(n140), .ZN(Z[7]) );
  AOI22_X1 U63 ( .A1(D[7]), .A2(n80), .B1(C[7]), .B2(n77), .ZN(n140) );
  NAND2_X1 U64 ( .A1(n143), .A2(n142), .ZN(Z[8]) );
  AOI22_X1 U65 ( .A1(D[8]), .A2(n80), .B1(C[8]), .B2(n77), .ZN(n142) );
  NAND2_X1 U66 ( .A1(n149), .A2(n148), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(D[9]), .A2(n80), .B1(C[9]), .B2(n77), .ZN(n148) );
  NAND2_X1 U68 ( .A1(n95), .A2(n94), .ZN(Z[15]) );
  AOI22_X1 U69 ( .A1(D[15]), .A2(n78), .B1(C[15]), .B2(n75), .ZN(n94) );
  NAND2_X1 U70 ( .A1(n97), .A2(n96), .ZN(Z[16]) );
  AOI22_X1 U71 ( .A1(D[16]), .A2(n78), .B1(C[16]), .B2(n75), .ZN(n96) );
  NAND2_X1 U72 ( .A1(n99), .A2(n98), .ZN(Z[17]) );
  AOI22_X1 U73 ( .A1(D[17]), .A2(n78), .B1(C[17]), .B2(n75), .ZN(n98) );
  NAND2_X1 U74 ( .A1(n101), .A2(n100), .ZN(Z[18]) );
  AOI22_X1 U75 ( .A1(D[18]), .A2(n78), .B1(C[18]), .B2(n75), .ZN(n100) );
  NAND2_X1 U76 ( .A1(n103), .A2(n102), .ZN(Z[19]) );
  AOI22_X1 U77 ( .A1(D[19]), .A2(n78), .B1(C[19]), .B2(n75), .ZN(n102) );
  NAND2_X1 U78 ( .A1(n107), .A2(n106), .ZN(Z[20]) );
  AOI22_X1 U79 ( .A1(D[20]), .A2(n79), .B1(C[20]), .B2(n76), .ZN(n106) );
  NAND2_X1 U80 ( .A1(n109), .A2(n108), .ZN(Z[21]) );
  AOI22_X1 U81 ( .A1(D[21]), .A2(n79), .B1(C[21]), .B2(n76), .ZN(n108) );
  NAND2_X1 U82 ( .A1(n111), .A2(n110), .ZN(Z[22]) );
  AOI22_X1 U83 ( .A1(D[22]), .A2(n79), .B1(C[22]), .B2(n76), .ZN(n110) );
  NAND2_X1 U84 ( .A1(n113), .A2(n112), .ZN(Z[23]) );
  AOI22_X1 U85 ( .A1(D[23]), .A2(n79), .B1(C[23]), .B2(n76), .ZN(n112) );
  NAND2_X1 U86 ( .A1(n115), .A2(n114), .ZN(Z[24]) );
  AOI22_X1 U87 ( .A1(D[24]), .A2(n79), .B1(C[24]), .B2(n76), .ZN(n114) );
  NAND2_X1 U88 ( .A1(n117), .A2(n116), .ZN(Z[25]) );
  AOI22_X1 U89 ( .A1(D[25]), .A2(n79), .B1(C[25]), .B2(n76), .ZN(n116) );
  NAND2_X1 U90 ( .A1(n119), .A2(n118), .ZN(Z[26]) );
  AOI22_X1 U91 ( .A1(D[26]), .A2(n79), .B1(C[26]), .B2(n76), .ZN(n118) );
  NAND2_X1 U92 ( .A1(n121), .A2(n120), .ZN(Z[27]) );
  AOI22_X1 U93 ( .A1(D[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n120) );
  NAND2_X1 U94 ( .A1(n123), .A2(n122), .ZN(Z[28]) );
  AOI22_X1 U95 ( .A1(D[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n122) );
  NAND2_X1 U96 ( .A1(n125), .A2(n124), .ZN(Z[29]) );
  AOI22_X1 U97 ( .A1(D[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n124) );
  NAND2_X1 U98 ( .A1(n129), .A2(n128), .ZN(Z[30]) );
  AOI22_X1 U99 ( .A1(D[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n128) );
  NAND2_X1 U100 ( .A1(n93), .A2(n92), .ZN(Z[14]) );
  AOI22_X1 U101 ( .A1(D[14]), .A2(n78), .B1(C[14]), .B2(n75), .ZN(n92) );
  NAND2_X1 U102 ( .A1(n105), .A2(n104), .ZN(Z[1]) );
  AOI22_X1 U103 ( .A1(D[1]), .A2(n78), .B1(C[1]), .B2(n75), .ZN(n104) );
  NAND2_X1 U104 ( .A1(n127), .A2(n126), .ZN(Z[2]) );
  AOI22_X1 U105 ( .A1(D[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n126) );
  NAND2_X1 U106 ( .A1(n85), .A2(n84), .ZN(Z[10]) );
  AOI22_X1 U107 ( .A1(D[10]), .A2(n78), .B1(C[10]), .B2(n75), .ZN(n84) );
  NAND2_X1 U108 ( .A1(n87), .A2(n86), .ZN(Z[11]) );
  AOI22_X1 U109 ( .A1(D[11]), .A2(n78), .B1(C[11]), .B2(n75), .ZN(n86) );
  NAND2_X1 U110 ( .A1(n89), .A2(n88), .ZN(Z[12]) );
  AOI22_X1 U111 ( .A1(D[12]), .A2(n78), .B1(C[12]), .B2(n75), .ZN(n88) );
  NAND2_X1 U112 ( .A1(n91), .A2(n90), .ZN(Z[13]) );
  AOI22_X1 U113 ( .A1(D[13]), .A2(n78), .B1(C[13]), .B2(n75), .ZN(n90) );
endmodule


module mux21_NBIT32_2 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  INV_X1 U12 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U13 ( .A1(A[31]), .A2(n4), .B1(B[31]), .B2(n7), .ZN(n103) );
  BUF_X1 U14 ( .A(S), .Z(n3) );
  BUF_X1 U15 ( .A(S), .Z(n2) );
  BUF_X1 U16 ( .A(S), .Z(n1) );
  INV_X1 U17 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U18 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U19 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U20 ( .A1(A[3]), .A2(n5), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U21 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U22 ( .A1(A[4]), .A2(n4), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U23 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U24 ( .A1(A[5]), .A2(n5), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U25 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U26 ( .A1(A[6]), .A2(n4), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U27 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U28 ( .A1(A[7]), .A2(n5), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U29 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U30 ( .A1(A[8]), .A2(n4), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U31 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U32 ( .A1(A[9]), .A2(n5), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U33 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U34 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U35 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U36 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U37 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U38 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U39 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U40 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U41 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U42 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U43 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U44 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U45 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U46 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U47 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U48 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U49 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U50 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U51 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U52 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U53 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U54 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U55 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U56 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U57 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U58 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U59 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U60 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U61 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U63 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U64 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U65 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U66 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U67 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U68 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U69 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U70 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U71 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U72 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U73 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U74 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U75 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U76 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U77 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U78 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
endmodule


module mux21_NBIT32_1 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n2) );
  BUF_X1 U14 ( .A(S), .Z(n1) );
  INV_X1 U15 ( .A(n79), .ZN(Z[0]) );
  AOI22_X1 U16 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(n13), .ZN(n79) );
  INV_X1 U17 ( .A(n90), .ZN(Z[1]) );
  AOI22_X1 U18 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(n10), .ZN(n90) );
  INV_X1 U19 ( .A(n101), .ZN(Z[2]) );
  AOI22_X1 U20 ( .A1(A[2]), .A2(n5), .B1(B[2]), .B2(n7), .ZN(n101) );
  INV_X1 U21 ( .A(n104), .ZN(Z[3]) );
  AOI22_X1 U22 ( .A1(A[3]), .A2(n4), .B1(B[3]), .B2(n7), .ZN(n104) );
  INV_X1 U23 ( .A(n105), .ZN(Z[4]) );
  AOI22_X1 U24 ( .A1(A[4]), .A2(n5), .B1(B[4]), .B2(n7), .ZN(n105) );
  INV_X1 U25 ( .A(n106), .ZN(Z[5]) );
  AOI22_X1 U26 ( .A1(A[5]), .A2(n4), .B1(B[5]), .B2(n6), .ZN(n106) );
  INV_X1 U27 ( .A(n107), .ZN(Z[6]) );
  AOI22_X1 U28 ( .A1(A[6]), .A2(n5), .B1(B[6]), .B2(n6), .ZN(n107) );
  INV_X1 U29 ( .A(n108), .ZN(Z[7]) );
  AOI22_X1 U30 ( .A1(A[7]), .A2(n4), .B1(B[7]), .B2(n6), .ZN(n108) );
  INV_X1 U31 ( .A(n109), .ZN(Z[8]) );
  AOI22_X1 U32 ( .A1(A[8]), .A2(n5), .B1(B[8]), .B2(n6), .ZN(n109) );
  INV_X1 U33 ( .A(n110), .ZN(Z[9]) );
  AOI22_X1 U34 ( .A1(A[9]), .A2(n4), .B1(n13), .B2(B[9]), .ZN(n110) );
  INV_X1 U35 ( .A(n80), .ZN(Z[10]) );
  AOI22_X1 U36 ( .A1(A[10]), .A2(n4), .B1(B[10]), .B2(n13), .ZN(n80) );
  INV_X1 U37 ( .A(n81), .ZN(Z[11]) );
  AOI22_X1 U38 ( .A1(A[11]), .A2(n4), .B1(B[11]), .B2(n13), .ZN(n81) );
  INV_X1 U39 ( .A(n82), .ZN(Z[12]) );
  AOI22_X1 U40 ( .A1(A[12]), .A2(n4), .B1(B[12]), .B2(n12), .ZN(n82) );
  INV_X1 U41 ( .A(n83), .ZN(Z[13]) );
  AOI22_X1 U42 ( .A1(A[13]), .A2(n4), .B1(B[13]), .B2(n12), .ZN(n83) );
  INV_X1 U43 ( .A(n84), .ZN(Z[14]) );
  AOI22_X1 U44 ( .A1(A[14]), .A2(n4), .B1(B[14]), .B2(n12), .ZN(n84) );
  INV_X1 U45 ( .A(n85), .ZN(Z[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n4), .B1(B[15]), .B2(n12), .ZN(n85) );
  INV_X1 U47 ( .A(n86), .ZN(Z[16]) );
  AOI22_X1 U48 ( .A1(A[16]), .A2(n4), .B1(B[16]), .B2(n11), .ZN(n86) );
  INV_X1 U49 ( .A(n87), .ZN(Z[17]) );
  AOI22_X1 U50 ( .A1(A[17]), .A2(n4), .B1(B[17]), .B2(n11), .ZN(n87) );
  INV_X1 U51 ( .A(n88), .ZN(Z[18]) );
  AOI22_X1 U52 ( .A1(A[18]), .A2(n4), .B1(B[18]), .B2(n11), .ZN(n88) );
  INV_X1 U53 ( .A(n89), .ZN(Z[19]) );
  AOI22_X1 U54 ( .A1(A[19]), .A2(n4), .B1(B[19]), .B2(n11), .ZN(n89) );
  INV_X1 U55 ( .A(n91), .ZN(Z[20]) );
  AOI22_X1 U56 ( .A1(A[20]), .A2(n5), .B1(B[20]), .B2(n10), .ZN(n91) );
  INV_X1 U57 ( .A(n92), .ZN(Z[21]) );
  AOI22_X1 U58 ( .A1(A[21]), .A2(n5), .B1(B[21]), .B2(n10), .ZN(n92) );
  INV_X1 U59 ( .A(n93), .ZN(Z[22]) );
  AOI22_X1 U60 ( .A1(A[22]), .A2(n5), .B1(B[22]), .B2(n9), .ZN(n93) );
  INV_X1 U61 ( .A(n94), .ZN(Z[23]) );
  AOI22_X1 U62 ( .A1(A[23]), .A2(n5), .B1(B[23]), .B2(n9), .ZN(n94) );
  INV_X1 U63 ( .A(n95), .ZN(Z[24]) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n5), .B1(B[24]), .B2(n9), .ZN(n95) );
  INV_X1 U65 ( .A(n96), .ZN(Z[25]) );
  AOI22_X1 U66 ( .A1(A[25]), .A2(n5), .B1(B[25]), .B2(n9), .ZN(n96) );
  INV_X1 U67 ( .A(n97), .ZN(Z[26]) );
  AOI22_X1 U68 ( .A1(A[26]), .A2(n5), .B1(B[26]), .B2(n8), .ZN(n97) );
  INV_X1 U69 ( .A(n98), .ZN(Z[27]) );
  AOI22_X1 U70 ( .A1(A[27]), .A2(n5), .B1(B[27]), .B2(n8), .ZN(n98) );
  INV_X1 U71 ( .A(n99), .ZN(Z[28]) );
  AOI22_X1 U72 ( .A1(A[28]), .A2(n5), .B1(B[28]), .B2(n8), .ZN(n99) );
  INV_X1 U73 ( .A(n100), .ZN(Z[29]) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n5), .B1(B[29]), .B2(n8), .ZN(n100) );
  INV_X1 U75 ( .A(n102), .ZN(Z[30]) );
  AOI22_X1 U76 ( .A1(A[30]), .A2(n5), .B1(B[30]), .B2(n10), .ZN(n102) );
  INV_X1 U77 ( .A(n103), .ZN(Z[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n5), .B1(B[31]), .B2(n7), .ZN(n103) );
endmodule


module ALU_NBIT32 ( OP1, OP2, ALU_OPC, ALU_RES );
  input [31:0] OP1;
  input [31:0] OP2;
  input [4:0] ALU_OPC;
  output [31:0] ALU_RES;
  wire   select_zero_sig, LOGIC_ARITH, LEFT_RIGHT, ADD_SUB, n78, n79, n80, n81,
         n82, n83, n84, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n85,
         n86, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31;
  wire   [1:0] select_type_sig;
  wire   [31:0] A_CMP;
  wire   [31:0] B_CMP;
  wire   [31:0] A_SHF;
  wire   [31:0] B_SHF;
  wire   [31:0] A_ADD;
  wire   [31:0] B_ADD;
  wire   [15:0] A_MUL;
  wire   [15:0] B_MUL;
  wire   [1:0] OPSel;
  wire   [31:0] LOGIC_RES;
  wire   [31:0] COMP_RES;
  wire   [31:0] SHIFT_RES;
  wire   [31:0] ADD_SUB_RES;
  wire   [31:0] MUL_RES;
  wire   [31:0] sig_intraMux;
  wire   [31:0] sig_ALU_RES;

  OAI22_X2 U227 ( .A1(n191), .A2(n35), .B1(n41), .B2(n68), .ZN(A_SHF[31]) );
  NOR2_X2 U257 ( .A1(n75), .A2(n26), .ZN(A_MUL[9]) );
  NOR2_X2 U258 ( .A1(n74), .A2(n26), .ZN(A_MUL[8]) );
  NOR2_X2 U259 ( .A1(n73), .A2(n26), .ZN(A_MUL[7]) );
  NOR2_X2 U260 ( .A1(n72), .A2(n26), .ZN(A_MUL[6]) );
  NOR2_X2 U261 ( .A1(n71), .A2(n25), .ZN(A_MUL[5]) );
  NOR2_X2 U262 ( .A1(n70), .A2(n25), .ZN(A_MUL[4]) );
  NOR2_X2 U263 ( .A1(n69), .A2(n25), .ZN(A_MUL[3]) );
  NOR2_X2 U264 ( .A1(n66), .A2(n25), .ZN(A_MUL[2]) );
  NOR2_X2 U265 ( .A1(n55), .A2(n25), .ZN(A_MUL[1]) );
  NOR2_X2 U267 ( .A1(n49), .A2(n25), .ZN(A_MUL[14]) );
  NOR2_X2 U268 ( .A1(n48), .A2(n25), .ZN(A_MUL[13]) );
  NOR2_X2 U269 ( .A1(n47), .A2(n25), .ZN(A_MUL[12]) );
  NOR2_X2 U270 ( .A1(n46), .A2(n25), .ZN(A_MUL[11]) );
  NOR2_X2 U271 ( .A1(n45), .A2(n25), .ZN(A_MUL[10]) );
  NOR2_X2 U272 ( .A1(n44), .A2(n25), .ZN(A_MUL[0]) );
  NAND3_X1 U427 ( .A1(n209), .A2(n208), .A3(n80), .ZN(n79) );
  NAND3_X1 U428 ( .A1(n43), .A2(n37), .A3(n34), .ZN(select_type_sig[1]) );
  NAND3_X1 U429 ( .A1(n84), .A2(n3), .A3(n34), .ZN(select_type_sig[0]) );
  NAND3_X1 U430 ( .A1(ALU_OPC[3]), .A2(n209), .A3(n156), .ZN(n84) );
  NAND3_X1 U431 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[3]), .A3(n156), .ZN(n158) );
  NAND3_X1 U432 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[1]), .A3(n162), .ZN(n82) );
  NAND3_X1 U434 ( .A1(n208), .A2(n206), .A3(ALU_OPC[4]), .ZN(n164) );
  OAI33_X1 U435 ( .A1(n208), .A2(n202), .A3(n209), .B1(n170), .B2(ALU_OPC[0]), 
        .B3(n207), .ZN(ADD_SUB) );
  NAND3_X1 U436 ( .A1(n206), .A2(n201), .A3(n208), .ZN(n170) );
  comparator_NBIT32 Comp ( .A(A_CMP), .B(B_CMP), .OPSel({n203, OPSel}), .RES({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, COMP_RES[0]}) );
  shifter_NBIT32 Shift ( .A(A_SHF), .B(B_SHF), .LOGIC_ARITH(LOGIC_ARITH), 
        .LEFT_RIGHT(LEFT_RIGHT), .RES(SHIFT_RES) );
  P4Adder_NBIT32 Add_Sub_unit ( .A(A_ADD), .B(B_ADD), .Cin(n2), .S(ADD_SUB_RES) );
  BOOTHMUL_numBit16 Booth_mul ( .A(A_MUL), .B(B_MUL), .P(MUL_RES) );
  mux41_NBIT32_1 Res_mux ( .A(ADD_SUB_RES), .B(LOGIC_RES), .C(SHIFT_RES), .D({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, COMP_RES[0]}), .S(
        select_type_sig), .Z(sig_intraMux) );
  mux21_NBIT32_2 Mul_mux ( .A(sig_intraMux), .B(MUL_RES), .S(n1), .Z(
        sig_ALU_RES) );
  mux21_NBIT32_1 Zeros_mux ( .A(sig_ALU_RES), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .S(select_zero_sig), .Z(ALU_RES) );
  OAI22_X1 U3 ( .A1(n194), .A2(n35), .B1(n40), .B2(n71), .ZN(A_SHF[5]) );
  OAI22_X1 U4 ( .A1(n195), .A2(n35), .B1(n40), .B2(n72), .ZN(A_SHF[6]) );
  OAI22_X1 U5 ( .A1(n185), .A2(n36), .B1(n41), .B2(n62), .ZN(A_SHF[26]) );
  OAI22_X1 U6 ( .A1(n186), .A2(n36), .B1(n41), .B2(n63), .ZN(A_SHF[27]) );
  AND3_X1 U7 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[2]), .A3(n163), .ZN(n1) );
  INV_X1 U8 ( .A(n199), .ZN(n2) );
  BUF_X1 U9 ( .A(n168), .Z(n13) );
  BUF_X1 U10 ( .A(n168), .Z(n14) );
  BUF_X1 U11 ( .A(n168), .Z(n15) );
  OAI22_X1 U12 ( .A1(n175), .A2(n37), .B1(n42), .B2(n52), .ZN(A_SHF[17]) );
  OAI22_X1 U13 ( .A1(n196), .A2(n35), .B1(n40), .B2(n73), .ZN(A_SHF[7]) );
  OAI22_X1 U14 ( .A1(n176), .A2(n37), .B1(n42), .B2(n53), .ZN(A_SHF[18]) );
  OAI22_X1 U15 ( .A1(n184), .A2(n36), .B1(n41), .B2(n61), .ZN(A_SHF[25]) );
  OAI22_X1 U16 ( .A1(n187), .A2(n36), .B1(n41), .B2(n64), .ZN(A_SHF[28]) );
  OAI22_X1 U17 ( .A1(n193), .A2(n36), .B1(n41), .B2(n70), .ZN(A_SHF[4]) );
  NOR2_X1 U18 ( .A1(n38), .A2(n192), .ZN(B_SHF[3]) );
  OAI22_X1 U19 ( .A1(n197), .A2(n35), .B1(n40), .B2(n74), .ZN(A_SHF[8]) );
  OAI22_X1 U20 ( .A1(n189), .A2(n35), .B1(n41), .B2(n66), .ZN(A_SHF[2]) );
  OAI22_X1 U21 ( .A1(n182), .A2(n36), .B1(n41), .B2(n59), .ZN(A_SHF[23]) );
  OAI22_X1 U22 ( .A1(n183), .A2(n36), .B1(n41), .B2(n60), .ZN(A_SHF[24]) );
  OAI22_X1 U23 ( .A1(n177), .A2(n36), .B1(n42), .B2(n54), .ZN(A_SHF[19]) );
  OAI22_X1 U24 ( .A1(n179), .A2(n36), .B1(n42), .B2(n56), .ZN(A_SHF[20]) );
  OAI22_X1 U25 ( .A1(n180), .A2(n36), .B1(n42), .B2(n57), .ZN(A_SHF[21]) );
  OAI22_X1 U26 ( .A1(n181), .A2(n36), .B1(n42), .B2(n58), .ZN(A_SHF[22]) );
  OAI22_X1 U27 ( .A1(n86), .A2(n37), .B1(n43), .B2(n47), .ZN(A_SHF[12]) );
  OAI22_X1 U28 ( .A1(n171), .A2(n37), .B1(n42), .B2(n48), .ZN(A_SHF[13]) );
  OAI22_X1 U29 ( .A1(n172), .A2(n37), .B1(n42), .B2(n49), .ZN(A_SHF[14]) );
  NOR2_X1 U30 ( .A1(n192), .A2(n26), .ZN(B_MUL[3]) );
  NOR2_X1 U31 ( .A1(n194), .A2(n26), .ZN(B_MUL[5]) );
  NOR2_X1 U32 ( .A1(n196), .A2(n26), .ZN(B_MUL[7]) );
  NOR2_X1 U33 ( .A1(n198), .A2(n26), .ZN(B_MUL[9]) );
  NOR2_X1 U34 ( .A1(n178), .A2(n26), .ZN(B_MUL[1]) );
  NOR2_X1 U35 ( .A1(n85), .A2(n26), .ZN(B_MUL[11]) );
  NOR2_X1 U36 ( .A1(n171), .A2(n26), .ZN(B_MUL[13]) );
  NOR2_X1 U37 ( .A1(n38), .A2(n198), .ZN(B_SHF[9]) );
  NOR2_X1 U38 ( .A1(n38), .A2(n197), .ZN(B_SHF[8]) );
  NOR2_X1 U39 ( .A1(n40), .A2(n77), .ZN(B_SHF[10]) );
  OAI22_X1 U40 ( .A1(n178), .A2(n36), .B1(n42), .B2(n55), .ZN(A_SHF[1]) );
  NOR2_X1 U41 ( .A1(n38), .A2(n189), .ZN(B_SHF[2]) );
  OAI22_X1 U42 ( .A1(n198), .A2(n35), .B1(n40), .B2(n75), .ZN(A_SHF[9]) );
  OAI22_X1 U43 ( .A1(n76), .A2(n35), .B1(n42), .B2(n44), .ZN(A_SHF[0]) );
  NOR2_X1 U44 ( .A1(n38), .A2(n196), .ZN(B_SHF[7]) );
  NOR2_X1 U45 ( .A1(n38), .A2(n195), .ZN(B_SHF[6]) );
  NOR2_X1 U46 ( .A1(n38), .A2(n194), .ZN(B_SHF[5]) );
  OAI22_X1 U47 ( .A1(n85), .A2(n37), .B1(n43), .B2(n46), .ZN(A_SHF[11]) );
  OAI22_X1 U48 ( .A1(n173), .A2(n37), .B1(n42), .B2(n50), .ZN(A_SHF[15]) );
  OAI22_X1 U49 ( .A1(n188), .A2(n35), .B1(n41), .B2(n65), .ZN(A_SHF[29]) );
  OAI22_X1 U50 ( .A1(n174), .A2(n37), .B1(n42), .B2(n51), .ZN(A_SHF[16]) );
  OAI22_X1 U51 ( .A1(n192), .A2(n35), .B1(n41), .B2(n69), .ZN(A_SHF[3]) );
  NOR2_X1 U52 ( .A1(n13), .A2(n44), .ZN(A_ADD[0]) );
  NOR2_X1 U53 ( .A1(n15), .A2(n70), .ZN(A_ADD[4]) );
  NOR2_X1 U54 ( .A1(n15), .A2(n74), .ZN(A_ADD[8]) );
  NOR2_X1 U55 ( .A1(n15), .A2(n71), .ZN(A_ADD[5]) );
  NOR2_X1 U56 ( .A1(n15), .A2(n75), .ZN(A_ADD[9]) );
  NOR2_X1 U57 ( .A1(n15), .A2(n72), .ZN(A_ADD[6]) );
  NOR2_X1 U58 ( .A1(n15), .A2(n69), .ZN(A_ADD[3]) );
  NOR2_X1 U59 ( .A1(n15), .A2(n73), .ZN(A_ADD[7]) );
  NOR2_X1 U60 ( .A1(n15), .A2(n68), .ZN(A_ADD[31]) );
  NOR2_X1 U61 ( .A1(n13), .A2(n47), .ZN(A_ADD[12]) );
  NOR2_X1 U62 ( .A1(n13), .A2(n51), .ZN(A_ADD[16]) );
  NOR2_X1 U63 ( .A1(n14), .A2(n60), .ZN(A_ADD[24]) );
  NOR2_X1 U64 ( .A1(n13), .A2(n55), .ZN(A_ADD[1]) );
  NOR2_X1 U65 ( .A1(n13), .A2(n48), .ZN(A_ADD[13]) );
  NOR2_X1 U66 ( .A1(n13), .A2(n52), .ZN(A_ADD[17]) );
  NOR2_X1 U67 ( .A1(n14), .A2(n61), .ZN(A_ADD[25]) );
  NOR2_X1 U68 ( .A1(n14), .A2(n66), .ZN(A_ADD[2]) );
  NOR2_X1 U69 ( .A1(n13), .A2(n45), .ZN(A_ADD[10]) );
  NOR2_X1 U70 ( .A1(n13), .A2(n49), .ZN(A_ADD[14]) );
  NOR2_X1 U71 ( .A1(n13), .A2(n53), .ZN(A_ADD[18]) );
  NOR2_X1 U72 ( .A1(n14), .A2(n62), .ZN(A_ADD[26]) );
  NOR2_X1 U73 ( .A1(n14), .A2(n58), .ZN(A_ADD[22]) );
  NOR2_X1 U74 ( .A1(n14), .A2(n57), .ZN(A_ADD[21]) );
  NOR2_X1 U75 ( .A1(n14), .A2(n56), .ZN(A_ADD[20]) );
  NOR2_X1 U76 ( .A1(n14), .A2(n67), .ZN(A_ADD[30]) );
  NOR2_X1 U77 ( .A1(n14), .A2(n65), .ZN(A_ADD[29]) );
  NOR2_X1 U78 ( .A1(n14), .A2(n64), .ZN(A_ADD[28]) );
  NOR2_X1 U79 ( .A1(n13), .A2(n46), .ZN(A_ADD[11]) );
  NOR2_X1 U80 ( .A1(n13), .A2(n50), .ZN(A_ADD[15]) );
  NOR2_X1 U81 ( .A1(n13), .A2(n54), .ZN(A_ADD[19]) );
  NOR2_X1 U82 ( .A1(n14), .A2(n59), .ZN(A_ADD[23]) );
  NOR2_X1 U83 ( .A1(n14), .A2(n63), .ZN(A_ADD[27]) );
  NOR2_X1 U84 ( .A1(n39), .A2(n178), .ZN(B_SHF[1]) );
  NOR2_X1 U85 ( .A1(n38), .A2(n187), .ZN(B_SHF[28]) );
  NOR2_X1 U86 ( .A1(n38), .A2(n186), .ZN(B_SHF[27]) );
  NOR2_X1 U87 ( .A1(n39), .A2(n185), .ZN(B_SHF[26]) );
  OAI22_X1 U88 ( .A1(n77), .A2(n37), .B1(n43), .B2(n45), .ZN(A_SHF[10]) );
  NOR2_X1 U89 ( .A1(n40), .A2(n85), .ZN(B_SHF[11]) );
  NOR2_X1 U90 ( .A1(n173), .A2(n26), .ZN(B_MUL[15]) );
  OAI22_X1 U91 ( .A1(n190), .A2(n35), .B1(n41), .B2(n67), .ZN(A_SHF[30]) );
  NOR2_X1 U92 ( .A1(n39), .A2(n176), .ZN(B_SHF[18]) );
  NOR2_X1 U93 ( .A1(n38), .A2(n188), .ZN(B_SHF[29]) );
  NOR2_X1 U94 ( .A1(n38), .A2(n190), .ZN(B_SHF[30]) );
  BUF_X1 U95 ( .A(n205), .Z(n7) );
  BUF_X1 U96 ( .A(n205), .Z(n8) );
  BUF_X1 U97 ( .A(n205), .Z(n9) );
  BUF_X1 U98 ( .A(n205), .Z(n11) );
  BUF_X1 U99 ( .A(n205), .Z(n10) );
  NOR2_X1 U100 ( .A1(n39), .A2(n184), .ZN(B_SHF[25]) );
  NOR2_X1 U101 ( .A1(n40), .A2(n76), .ZN(B_SHF[0]) );
  NOR2_X1 U102 ( .A1(n39), .A2(n174), .ZN(B_SHF[16]) );
  NOR2_X1 U103 ( .A1(n39), .A2(n175), .ZN(B_SHF[17]) );
  NOR2_X1 U104 ( .A1(n40), .A2(n173), .ZN(B_SHF[15]) );
  NOR2_X1 U105 ( .A1(n50), .A2(n25), .ZN(A_MUL[15]) );
  NOR2_X1 U106 ( .A1(n189), .A2(n26), .ZN(B_MUL[2]) );
  NOR2_X1 U107 ( .A1(n193), .A2(n25), .ZN(B_MUL[4]) );
  NOR2_X1 U108 ( .A1(n195), .A2(n26), .ZN(B_MUL[6]) );
  NOR2_X1 U109 ( .A1(n197), .A2(n25), .ZN(B_MUL[8]) );
  NOR2_X1 U110 ( .A1(n76), .A2(n26), .ZN(B_MUL[0]) );
  NOR2_X1 U111 ( .A1(n77), .A2(n26), .ZN(B_MUL[10]) );
  NOR2_X1 U112 ( .A1(n86), .A2(n26), .ZN(B_MUL[12]) );
  NOR2_X1 U113 ( .A1(n172), .A2(n26), .ZN(B_MUL[14]) );
  BUF_X1 U114 ( .A(n199), .Z(n5) );
  BUF_X1 U115 ( .A(n199), .Z(n4) );
  OAI21_X1 U116 ( .B1(n43), .B2(n193), .A(n37), .ZN(B_SHF[4]) );
  BUF_X1 U117 ( .A(n199), .Z(n6) );
  NOR2_X1 U118 ( .A1(n39), .A2(n183), .ZN(B_SHF[24]) );
  NOR2_X1 U119 ( .A1(n39), .A2(n182), .ZN(B_SHF[23]) );
  NOR2_X1 U120 ( .A1(n39), .A2(n181), .ZN(B_SHF[22]) );
  NOR2_X1 U121 ( .A1(n30), .A2(n67), .ZN(A_CMP[30]) );
  OAI22_X1 U122 ( .A1(n99), .A2(n194), .B1(n100), .B2(n71), .ZN(LOGIC_RES[5])
         );
  OAI22_X1 U123 ( .A1(n97), .A2(n195), .B1(n98), .B2(n72), .ZN(LOGIC_RES[6])
         );
  OAI22_X1 U124 ( .A1(n95), .A2(n196), .B1(n96), .B2(n73), .ZN(LOGIC_RES[7])
         );
  OAI22_X1 U125 ( .A1(n90), .A2(n198), .B1(n91), .B2(n75), .ZN(LOGIC_RES[9])
         );
  OAI22_X1 U126 ( .A1(n105), .A2(n191), .B1(n106), .B2(n68), .ZN(LOGIC_RES[31]) );
  NOR2_X1 U127 ( .A1(n29), .A2(n55), .ZN(A_CMP[1]) );
  OAI22_X1 U128 ( .A1(n151), .A2(n77), .B1(n152), .B2(n45), .ZN(LOGIC_RES[10])
         );
  OAI22_X1 U129 ( .A1(n149), .A2(n85), .B1(n150), .B2(n46), .ZN(LOGIC_RES[11])
         );
  OAI22_X1 U130 ( .A1(n145), .A2(n171), .B1(n146), .B2(n48), .ZN(LOGIC_RES[13]) );
  OAI22_X1 U131 ( .A1(n143), .A2(n172), .B1(n144), .B2(n49), .ZN(LOGIC_RES[14]) );
  OAI22_X1 U132 ( .A1(n141), .A2(n173), .B1(n142), .B2(n50), .ZN(LOGIC_RES[15]) );
  OAI22_X1 U133 ( .A1(n137), .A2(n175), .B1(n138), .B2(n52), .ZN(LOGIC_RES[17]) );
  OAI22_X1 U134 ( .A1(n135), .A2(n176), .B1(n136), .B2(n53), .ZN(LOGIC_RES[18]) );
  OAI22_X1 U135 ( .A1(n133), .A2(n177), .B1(n134), .B2(n54), .ZN(LOGIC_RES[19]) );
  OAI22_X1 U136 ( .A1(n127), .A2(n180), .B1(n128), .B2(n57), .ZN(LOGIC_RES[21]) );
  OAI22_X1 U137 ( .A1(n125), .A2(n181), .B1(n126), .B2(n58), .ZN(LOGIC_RES[22]) );
  OAI22_X1 U138 ( .A1(n123), .A2(n182), .B1(n124), .B2(n59), .ZN(LOGIC_RES[23]) );
  OAI22_X1 U139 ( .A1(n119), .A2(n184), .B1(n120), .B2(n61), .ZN(LOGIC_RES[25]) );
  OAI22_X1 U140 ( .A1(n117), .A2(n185), .B1(n118), .B2(n62), .ZN(LOGIC_RES[26]) );
  OAI22_X1 U141 ( .A1(n115), .A2(n186), .B1(n116), .B2(n63), .ZN(LOGIC_RES[27]) );
  OAI22_X1 U142 ( .A1(n111), .A2(n188), .B1(n112), .B2(n65), .ZN(LOGIC_RES[29]) );
  OAI22_X1 U143 ( .A1(n107), .A2(n190), .B1(n108), .B2(n67), .ZN(LOGIC_RES[30]) );
  NOR2_X1 U144 ( .A1(n39), .A2(n177), .ZN(B_SHF[19]) );
  NOR2_X1 U145 ( .A1(n39), .A2(n180), .ZN(B_SHF[21]) );
  NOR2_X1 U146 ( .A1(n40), .A2(n171), .ZN(B_SHF[13]) );
  NOR2_X1 U147 ( .A1(n39), .A2(n179), .ZN(B_SHF[20]) );
  NOR2_X1 U148 ( .A1(n40), .A2(n172), .ZN(B_SHF[14]) );
  NOR2_X1 U149 ( .A1(n40), .A2(n86), .ZN(B_SHF[12]) );
  NOR2_X1 U150 ( .A1(n34), .A2(n196), .ZN(B_CMP[7]) );
  NOR2_X1 U151 ( .A1(n34), .A2(n198), .ZN(B_CMP[9]) );
  AOI21_X1 U152 ( .B1(n9), .B2(n194), .A(n21), .ZN(n100) );
  AOI21_X1 U153 ( .B1(n9), .B2(n195), .A(n21), .ZN(n98) );
  AOI21_X1 U154 ( .B1(n9), .B2(n197), .A(n21), .ZN(n94) );
  AOI21_X1 U155 ( .B1(n11), .B2(n178), .A(n23), .ZN(n132) );
  AOI21_X1 U156 ( .B1(n10), .B2(n189), .A(n22), .ZN(n110) );
  AOI21_X1 U157 ( .B1(n10), .B2(n192), .A(n22), .ZN(n104) );
  AOI21_X1 U158 ( .B1(n10), .B2(n193), .A(n22), .ZN(n102) );
  AOI21_X1 U159 ( .B1(n10), .B2(n196), .A(n22), .ZN(n96) );
  AOI21_X1 U160 ( .B1(n10), .B2(n198), .A(n22), .ZN(n91) );
  AOI21_X1 U161 ( .B1(n11), .B2(n172), .A(n23), .ZN(n144) );
  AOI21_X1 U162 ( .B1(n11), .B2(n173), .A(n23), .ZN(n142) );
  AOI21_X1 U163 ( .B1(n11), .B2(n174), .A(n23), .ZN(n140) );
  AOI21_X1 U164 ( .B1(n11), .B2(n175), .A(n23), .ZN(n138) );
  AOI21_X1 U165 ( .B1(n11), .B2(n176), .A(n23), .ZN(n136) );
  AOI21_X1 U166 ( .B1(n11), .B2(n177), .A(n23), .ZN(n134) );
  AOI21_X1 U167 ( .B1(n11), .B2(n179), .A(n23), .ZN(n130) );
  AOI21_X1 U168 ( .B1(n11), .B2(n180), .A(n23), .ZN(n128) );
  AOI21_X1 U169 ( .B1(n11), .B2(n181), .A(n23), .ZN(n126) );
  AOI21_X1 U170 ( .B1(n11), .B2(n182), .A(n23), .ZN(n124) );
  AOI21_X1 U171 ( .B1(n11), .B2(n183), .A(n22), .ZN(n122) );
  AOI21_X1 U172 ( .B1(n10), .B2(n184), .A(n22), .ZN(n120) );
  AOI21_X1 U173 ( .B1(n10), .B2(n185), .A(n22), .ZN(n118) );
  AOI21_X1 U174 ( .B1(n10), .B2(n186), .A(n22), .ZN(n116) );
  AOI21_X1 U175 ( .B1(n10), .B2(n187), .A(n22), .ZN(n114) );
  AOI21_X1 U176 ( .B1(n10), .B2(n188), .A(n22), .ZN(n112) );
  AOI21_X1 U177 ( .B1(n10), .B2(n190), .A(n22), .ZN(n108) );
  AOI21_X1 U178 ( .B1(n10), .B2(n191), .A(n22), .ZN(n106) );
  AOI21_X1 U179 ( .B1(n12), .B2(n77), .A(n24), .ZN(n152) );
  AOI21_X1 U180 ( .B1(n12), .B2(n85), .A(n24), .ZN(n150) );
  AOI21_X1 U181 ( .B1(n12), .B2(n86), .A(n23), .ZN(n148) );
  AOI21_X1 U182 ( .B1(n12), .B2(n171), .A(n23), .ZN(n146) );
  NOR2_X1 U183 ( .A1(n34), .A2(n197), .ZN(B_CMP[8]) );
  NOR2_X1 U184 ( .A1(n34), .A2(n195), .ZN(B_CMP[6]) );
  NOR2_X1 U185 ( .A1(n33), .A2(n190), .ZN(B_CMP[30]) );
  NOR2_X1 U186 ( .A1(n31), .A2(n76), .ZN(B_CMP[0]) );
  NOR2_X1 U187 ( .A1(n33), .A2(n192), .ZN(B_CMP[3]) );
  NOR2_X1 U188 ( .A1(n33), .A2(n194), .ZN(B_CMP[5]) );
  NOR2_X1 U189 ( .A1(n31), .A2(n85), .ZN(B_CMP[11]) );
  NOR2_X1 U190 ( .A1(n32), .A2(n171), .ZN(B_CMP[13]) );
  NOR2_X1 U191 ( .A1(n32), .A2(n173), .ZN(B_CMP[15]) );
  NOR2_X1 U192 ( .A1(n32), .A2(n175), .ZN(B_CMP[17]) );
  NOR2_X1 U193 ( .A1(n32), .A2(n177), .ZN(B_CMP[19]) );
  NOR2_X1 U194 ( .A1(n32), .A2(n180), .ZN(B_CMP[21]) );
  NOR2_X1 U195 ( .A1(n32), .A2(n182), .ZN(B_CMP[23]) );
  NOR2_X1 U196 ( .A1(n33), .A2(n184), .ZN(B_CMP[25]) );
  NOR2_X1 U197 ( .A1(n33), .A2(n186), .ZN(B_CMP[27]) );
  NOR2_X1 U198 ( .A1(n33), .A2(n188), .ZN(B_CMP[29]) );
  NOR2_X1 U199 ( .A1(n31), .A2(n68), .ZN(A_CMP[31]) );
  NOR2_X1 U200 ( .A1(n33), .A2(n193), .ZN(B_CMP[4]) );
  NOR2_X1 U201 ( .A1(n31), .A2(n86), .ZN(B_CMP[12]) );
  NOR2_X1 U202 ( .A1(n32), .A2(n174), .ZN(B_CMP[16]) );
  NOR2_X1 U203 ( .A1(n32), .A2(n179), .ZN(B_CMP[20]) );
  NOR2_X1 U204 ( .A1(n33), .A2(n183), .ZN(B_CMP[24]) );
  NOR2_X1 U205 ( .A1(n33), .A2(n187), .ZN(B_CMP[28]) );
  NOR2_X1 U206 ( .A1(n33), .A2(n189), .ZN(B_CMP[2]) );
  NOR2_X1 U207 ( .A1(n31), .A2(n77), .ZN(B_CMP[10]) );
  NOR2_X1 U208 ( .A1(n32), .A2(n172), .ZN(B_CMP[14]) );
  NOR2_X1 U209 ( .A1(n32), .A2(n176), .ZN(B_CMP[18]) );
  NOR2_X1 U210 ( .A1(n32), .A2(n181), .ZN(B_CMP[22]) );
  NOR2_X1 U211 ( .A1(n33), .A2(n185), .ZN(B_CMP[26]) );
  AND2_X1 U212 ( .A1(n18), .A2(n6), .ZN(n168) );
  NOR2_X1 U213 ( .A1(n38), .A2(n191), .ZN(B_SHF[31]) );
  NOR2_X1 U214 ( .A1(n32), .A2(n178), .ZN(B_CMP[1]) );
  NOR2_X1 U215 ( .A1(n29), .A2(n44), .ZN(A_CMP[0]) );
  NOR2_X1 U216 ( .A1(n31), .A2(n69), .ZN(A_CMP[3]) );
  NOR2_X1 U217 ( .A1(n31), .A2(n71), .ZN(A_CMP[5]) );
  NOR2_X1 U218 ( .A1(n31), .A2(n73), .ZN(A_CMP[7]) );
  NOR2_X1 U219 ( .A1(n31), .A2(n75), .ZN(A_CMP[9]) );
  NOR2_X1 U220 ( .A1(n29), .A2(n46), .ZN(A_CMP[11]) );
  NOR2_X1 U221 ( .A1(n29), .A2(n48), .ZN(A_CMP[13]) );
  NOR2_X1 U222 ( .A1(n29), .A2(n50), .ZN(A_CMP[15]) );
  NOR2_X1 U223 ( .A1(n33), .A2(n191), .ZN(B_CMP[31]) );
  NOR2_X1 U224 ( .A1(n29), .A2(n52), .ZN(A_CMP[17]) );
  NOR2_X1 U225 ( .A1(n29), .A2(n54), .ZN(A_CMP[19]) );
  NOR2_X1 U226 ( .A1(n30), .A2(n57), .ZN(A_CMP[21]) );
  NOR2_X1 U228 ( .A1(n30), .A2(n59), .ZN(A_CMP[23]) );
  NOR2_X1 U229 ( .A1(n30), .A2(n61), .ZN(A_CMP[25]) );
  NOR2_X1 U230 ( .A1(n30), .A2(n63), .ZN(A_CMP[27]) );
  NOR2_X1 U231 ( .A1(n30), .A2(n65), .ZN(A_CMP[29]) );
  NOR2_X1 U232 ( .A1(n31), .A2(n70), .ZN(A_CMP[4]) );
  NOR2_X1 U233 ( .A1(n31), .A2(n74), .ZN(A_CMP[8]) );
  NOR2_X1 U234 ( .A1(n29), .A2(n47), .ZN(A_CMP[12]) );
  NOR2_X1 U235 ( .A1(n30), .A2(n66), .ZN(A_CMP[2]) );
  NOR2_X1 U236 ( .A1(n31), .A2(n72), .ZN(A_CMP[6]) );
  NOR2_X1 U237 ( .A1(n29), .A2(n45), .ZN(A_CMP[10]) );
  NOR2_X1 U238 ( .A1(n29), .A2(n49), .ZN(A_CMP[14]) );
  NOR2_X1 U239 ( .A1(n29), .A2(n51), .ZN(A_CMP[16]) );
  NOR2_X1 U240 ( .A1(n30), .A2(n56), .ZN(A_CMP[20]) );
  NOR2_X1 U241 ( .A1(n30), .A2(n60), .ZN(A_CMP[24]) );
  NOR2_X1 U242 ( .A1(n30), .A2(n64), .ZN(A_CMP[28]) );
  NOR2_X1 U243 ( .A1(n29), .A2(n53), .ZN(A_CMP[18]) );
  NOR2_X1 U244 ( .A1(n30), .A2(n58), .ZN(A_CMP[22]) );
  NOR2_X1 U245 ( .A1(n30), .A2(n62), .ZN(A_CMP[26]) );
  OAI22_X1 U246 ( .A1(OP2[0]), .A2(n6), .B1(n76), .B2(n18), .ZN(B_ADD[0]) );
  OAI22_X1 U247 ( .A1(OP2[4]), .A2(n4), .B1(n193), .B2(n16), .ZN(B_ADD[4]) );
  OAI22_X1 U248 ( .A1(OP2[8]), .A2(n4), .B1(n197), .B2(n16), .ZN(B_ADD[8]) );
  OAI22_X1 U249 ( .A1(OP2[12]), .A2(n6), .B1(n86), .B2(n18), .ZN(B_ADD[12]) );
  OAI22_X1 U250 ( .A1(OP2[16]), .A2(n6), .B1(n174), .B2(n18), .ZN(B_ADD[16])
         );
  OAI22_X1 U251 ( .A1(OP2[24]), .A2(n5), .B1(n183), .B2(n17), .ZN(B_ADD[24])
         );
  OAI22_X1 U252 ( .A1(OP2[5]), .A2(n4), .B1(n194), .B2(n16), .ZN(B_ADD[5]) );
  OAI22_X1 U253 ( .A1(OP2[1]), .A2(n5), .B1(n178), .B2(n17), .ZN(B_ADD[1]) );
  OAI22_X1 U254 ( .A1(OP2[9]), .A2(n4), .B1(n198), .B2(n16), .ZN(B_ADD[9]) );
  OAI22_X1 U255 ( .A1(OP2[13]), .A2(n6), .B1(n171), .B2(n18), .ZN(B_ADD[13])
         );
  OAI22_X1 U256 ( .A1(OP2[17]), .A2(n5), .B1(n175), .B2(n17), .ZN(B_ADD[17])
         );
  OAI22_X1 U266 ( .A1(OP2[25]), .A2(n5), .B1(n184), .B2(n17), .ZN(B_ADD[25])
         );
  OAI22_X1 U273 ( .A1(OP2[2]), .A2(n4), .B1(n189), .B2(n16), .ZN(B_ADD[2]) );
  OAI22_X1 U274 ( .A1(OP2[6]), .A2(n4), .B1(n195), .B2(n16), .ZN(B_ADD[6]) );
  OAI22_X1 U275 ( .A1(OP2[10]), .A2(n6), .B1(n77), .B2(n18), .ZN(B_ADD[10]) );
  OAI22_X1 U276 ( .A1(OP2[14]), .A2(n6), .B1(n172), .B2(n18), .ZN(B_ADD[14])
         );
  OAI22_X1 U277 ( .A1(OP2[18]), .A2(n5), .B1(n176), .B2(n17), .ZN(B_ADD[18])
         );
  OAI22_X1 U278 ( .A1(OP2[26]), .A2(n5), .B1(n185), .B2(n17), .ZN(B_ADD[26])
         );
  OAI22_X1 U279 ( .A1(OP2[22]), .A2(n5), .B1(n181), .B2(n17), .ZN(B_ADD[22])
         );
  OAI22_X1 U280 ( .A1(OP2[21]), .A2(n5), .B1(n180), .B2(n17), .ZN(B_ADD[21])
         );
  OAI22_X1 U281 ( .A1(OP2[20]), .A2(n5), .B1(n179), .B2(n17), .ZN(B_ADD[20])
         );
  OAI22_X1 U282 ( .A1(OP2[30]), .A2(n4), .B1(n190), .B2(n16), .ZN(B_ADD[30])
         );
  OAI22_X1 U283 ( .A1(OP2[29]), .A2(n4), .B1(n188), .B2(n16), .ZN(B_ADD[29])
         );
  OAI22_X1 U284 ( .A1(OP2[28]), .A2(n4), .B1(n187), .B2(n16), .ZN(B_ADD[28])
         );
  OAI22_X1 U285 ( .A1(OP2[3]), .A2(n4), .B1(n192), .B2(n16), .ZN(B_ADD[3]) );
  OAI22_X1 U286 ( .A1(OP2[7]), .A2(n4), .B1(n196), .B2(n16), .ZN(B_ADD[7]) );
  OAI22_X1 U287 ( .A1(OP2[11]), .A2(n6), .B1(n85), .B2(n18), .ZN(B_ADD[11]) );
  OAI22_X1 U288 ( .A1(OP2[15]), .A2(n6), .B1(n173), .B2(n18), .ZN(B_ADD[15])
         );
  OAI22_X1 U289 ( .A1(OP2[19]), .A2(n5), .B1(n177), .B2(n17), .ZN(B_ADD[19])
         );
  OAI22_X1 U290 ( .A1(OP2[23]), .A2(n5), .B1(n182), .B2(n17), .ZN(B_ADD[23])
         );
  OAI22_X1 U291 ( .A1(OP2[27]), .A2(n5), .B1(n186), .B2(n17), .ZN(B_ADD[27])
         );
  OAI22_X1 U292 ( .A1(OP2[31]), .A2(n4), .B1(n191), .B2(n16), .ZN(B_ADD[31])
         );
  INV_X1 U293 ( .A(n1), .ZN(n26) );
  INV_X1 U294 ( .A(n1), .ZN(n25) );
  INV_X1 U295 ( .A(n3), .ZN(n27) );
  INV_X1 U296 ( .A(n3), .ZN(n28) );
  INV_X1 U297 ( .A(ADD_SUB), .ZN(n199) );
  AOI221_X1 U298 ( .B1(OP1[10]), .B2(n27), .C1(n7), .C2(n45), .A(n19), .ZN(
        n151) );
  AOI221_X1 U299 ( .B1(OP1[11]), .B2(n28), .C1(n7), .C2(n46), .A(n19), .ZN(
        n149) );
  AOI221_X1 U300 ( .B1(OP1[12]), .B2(n27), .C1(n7), .C2(n47), .A(n19), .ZN(
        n147) );
  AOI221_X1 U301 ( .B1(OP1[13]), .B2(n28), .C1(n7), .C2(n48), .A(n19), .ZN(
        n145) );
  AOI221_X1 U302 ( .B1(OP1[14]), .B2(n27), .C1(n7), .C2(n49), .A(n19), .ZN(
        n143) );
  AOI221_X1 U303 ( .B1(OP1[15]), .B2(n28), .C1(n7), .C2(n50), .A(n19), .ZN(
        n141) );
  AOI221_X1 U304 ( .B1(OP1[16]), .B2(n27), .C1(n7), .C2(n51), .A(n19), .ZN(
        n139) );
  AOI221_X1 U305 ( .B1(OP1[1]), .B2(n28), .C1(n8), .C2(n55), .A(n20), .ZN(n131) );
  AOI221_X1 U306 ( .B1(OP1[2]), .B2(n27), .C1(n9), .C2(n66), .A(n21), .ZN(n109) );
  AOI221_X1 U307 ( .B1(OP1[3]), .B2(n27), .C1(n8), .C2(n69), .A(n20), .ZN(n103) );
  AOI221_X1 U308 ( .B1(OP1[4]), .B2(n27), .C1(n8), .C2(n70), .A(n20), .ZN(n101) );
  AOI221_X1 U309 ( .B1(OP1[5]), .B2(n27), .C1(n8), .C2(n71), .A(n20), .ZN(n99)
         );
  AOI221_X1 U310 ( .B1(OP1[6]), .B2(n27), .C1(n7), .C2(n72), .A(n19), .ZN(n97)
         );
  AOI221_X1 U311 ( .B1(OP1[7]), .B2(n27), .C1(n7), .C2(n73), .A(n19), .ZN(n95)
         );
  AOI221_X1 U312 ( .B1(OP1[8]), .B2(n27), .C1(n7), .C2(n74), .A(n19), .ZN(n93)
         );
  AOI221_X1 U313 ( .B1(OP1[17]), .B2(n28), .C1(n8), .C2(n52), .A(n20), .ZN(
        n137) );
  AOI221_X1 U314 ( .B1(OP1[18]), .B2(n28), .C1(n8), .C2(n53), .A(n20), .ZN(
        n135) );
  AOI221_X1 U315 ( .B1(OP1[19]), .B2(n28), .C1(n8), .C2(n54), .A(n20), .ZN(
        n133) );
  AOI221_X1 U316 ( .B1(OP1[20]), .B2(n28), .C1(n8), .C2(n56), .A(n20), .ZN(
        n129) );
  AOI221_X1 U317 ( .B1(OP1[21]), .B2(n28), .C1(n8), .C2(n57), .A(n20), .ZN(
        n127) );
  AOI221_X1 U318 ( .B1(OP1[22]), .B2(n28), .C1(n8), .C2(n58), .A(n20), .ZN(
        n125) );
  AOI221_X1 U319 ( .B1(OP1[23]), .B2(n28), .C1(n8), .C2(n59), .A(n20), .ZN(
        n123) );
  AOI221_X1 U320 ( .B1(OP1[24]), .B2(n28), .C1(n9), .C2(n60), .A(n21), .ZN(
        n121) );
  AOI221_X1 U321 ( .B1(OP1[25]), .B2(n28), .C1(n9), .C2(n61), .A(n21), .ZN(
        n119) );
  AOI221_X1 U322 ( .B1(OP1[26]), .B2(n28), .C1(n8), .C2(n62), .A(n20), .ZN(
        n117) );
  AOI221_X1 U323 ( .B1(OP1[27]), .B2(n28), .C1(n9), .C2(n63), .A(n21), .ZN(
        n115) );
  AOI221_X1 U324 ( .B1(OP1[28]), .B2(n27), .C1(n9), .C2(n64), .A(n21), .ZN(
        n113) );
  AOI221_X1 U325 ( .B1(OP1[29]), .B2(n27), .C1(n9), .C2(n65), .A(n21), .ZN(
        n111) );
  AOI221_X1 U326 ( .B1(OP1[30]), .B2(n27), .C1(n9), .C2(n67), .A(n21), .ZN(
        n107) );
  AOI221_X1 U327 ( .B1(OP1[31]), .B2(n27), .C1(n9), .C2(n68), .A(n21), .ZN(
        n105) );
  AOI221_X1 U328 ( .B1(n27), .B2(OP1[9]), .C1(n7), .C2(n75), .A(n19), .ZN(n90)
         );
  BUF_X1 U329 ( .A(n81), .Z(n39) );
  BUF_X1 U330 ( .A(n81), .Z(n40) );
  BUF_X1 U331 ( .A(n81), .Z(n41) );
  BUF_X1 U332 ( .A(n81), .Z(n42) );
  INV_X1 U333 ( .A(OP2[0]), .ZN(n76) );
  INV_X1 U334 ( .A(OP2[1]), .ZN(n178) );
  INV_X1 U335 ( .A(OP2[2]), .ZN(n189) );
  INV_X1 U336 ( .A(OP2[3]), .ZN(n192) );
  INV_X1 U337 ( .A(OP2[5]), .ZN(n194) );
  INV_X1 U338 ( .A(OP2[6]), .ZN(n195) );
  INV_X1 U339 ( .A(OP2[7]), .ZN(n196) );
  INV_X1 U340 ( .A(OP2[8]), .ZN(n197) );
  INV_X1 U341 ( .A(OP2[9]), .ZN(n198) );
  INV_X1 U342 ( .A(OP2[10]), .ZN(n77) );
  INV_X1 U343 ( .A(OP2[11]), .ZN(n85) );
  INV_X1 U344 ( .A(OP2[12]), .ZN(n86) );
  INV_X1 U345 ( .A(OP2[13]), .ZN(n171) );
  INV_X1 U346 ( .A(OP2[14]), .ZN(n172) );
  INV_X1 U347 ( .A(OP2[15]), .ZN(n173) );
  INV_X1 U348 ( .A(OP2[4]), .ZN(n193) );
  BUF_X1 U349 ( .A(n92), .Z(n19) );
  BUF_X1 U350 ( .A(n92), .Z(n20) );
  OAI22_X1 U351 ( .A1(n153), .A2(n76), .B1(n154), .B2(n44), .ZN(LOGIC_RES[0])
         );
  AOI21_X1 U352 ( .B1(n9), .B2(n76), .A(n21), .ZN(n154) );
  AOI221_X1 U353 ( .B1(OP1[0]), .B2(n28), .C1(n7), .C2(n44), .A(n19), .ZN(n153) );
  BUF_X1 U354 ( .A(n92), .Z(n23) );
  BUF_X1 U355 ( .A(n92), .Z(n22) );
  BUF_X1 U356 ( .A(n82), .Z(n35) );
  BUF_X1 U357 ( .A(n82), .Z(n36) );
  BUF_X1 U358 ( .A(n92), .Z(n21) );
  BUF_X1 U359 ( .A(n159), .Z(n17) );
  BUF_X1 U360 ( .A(n159), .Z(n16) );
  BUF_X1 U361 ( .A(n83), .Z(n33) );
  BUF_X1 U362 ( .A(n83), .Z(n31) );
  BUF_X1 U363 ( .A(n83), .Z(n29) );
  BUF_X1 U364 ( .A(n83), .Z(n32) );
  BUF_X1 U365 ( .A(n83), .Z(n30) );
  BUF_X1 U366 ( .A(n81), .Z(n38) );
  INV_X1 U367 ( .A(OP1[0]), .ZN(n44) );
  INV_X1 U368 ( .A(OP1[1]), .ZN(n55) );
  INV_X1 U369 ( .A(OP1[2]), .ZN(n66) );
  INV_X1 U370 ( .A(OP1[3]), .ZN(n69) );
  INV_X1 U371 ( .A(OP1[4]), .ZN(n70) );
  INV_X1 U372 ( .A(OP1[5]), .ZN(n71) );
  INV_X1 U373 ( .A(OP1[6]), .ZN(n72) );
  INV_X1 U374 ( .A(OP1[7]), .ZN(n73) );
  INV_X1 U375 ( .A(OP1[8]), .ZN(n74) );
  INV_X1 U376 ( .A(OP1[9]), .ZN(n75) );
  INV_X1 U377 ( .A(OP1[10]), .ZN(n45) );
  INV_X1 U378 ( .A(OP1[11]), .ZN(n46) );
  INV_X1 U379 ( .A(OP1[12]), .ZN(n47) );
  INV_X1 U380 ( .A(OP1[13]), .ZN(n48) );
  INV_X1 U381 ( .A(OP1[14]), .ZN(n49) );
  INV_X1 U382 ( .A(OP1[15]), .ZN(n50) );
  BUF_X1 U383 ( .A(n159), .Z(n18) );
  INV_X1 U384 ( .A(OP2[16]), .ZN(n174) );
  INV_X1 U385 ( .A(OP2[17]), .ZN(n175) );
  INV_X1 U386 ( .A(OP2[18]), .ZN(n176) );
  INV_X1 U387 ( .A(OP2[19]), .ZN(n177) );
  INV_X1 U388 ( .A(OP2[20]), .ZN(n179) );
  INV_X1 U389 ( .A(OP2[21]), .ZN(n180) );
  INV_X1 U390 ( .A(OP2[22]), .ZN(n181) );
  INV_X1 U391 ( .A(OP2[23]), .ZN(n182) );
  INV_X1 U392 ( .A(OP2[24]), .ZN(n183) );
  INV_X1 U393 ( .A(OP2[25]), .ZN(n184) );
  INV_X1 U394 ( .A(OP2[26]), .ZN(n185) );
  INV_X1 U395 ( .A(OP2[27]), .ZN(n186) );
  INV_X1 U396 ( .A(OP2[28]), .ZN(n187) );
  INV_X1 U397 ( .A(OP2[29]), .ZN(n188) );
  INV_X1 U398 ( .A(OP2[30]), .ZN(n190) );
  INV_X1 U399 ( .A(OP2[31]), .ZN(n191) );
  BUF_X1 U400 ( .A(n82), .Z(n37) );
  NAND2_X1 U401 ( .A1(n88), .A2(n89), .ZN(OPSel[0]) );
  OAI22_X1 U402 ( .A1(n103), .A2(n192), .B1(n104), .B2(n69), .ZN(LOGIC_RES[3])
         );
  OAI22_X1 U403 ( .A1(n101), .A2(n193), .B1(n102), .B2(n70), .ZN(LOGIC_RES[4])
         );
  OAI22_X1 U404 ( .A1(n93), .A2(n197), .B1(n94), .B2(n74), .ZN(LOGIC_RES[8])
         );
  OAI22_X1 U405 ( .A1(n131), .A2(n178), .B1(n132), .B2(n55), .ZN(LOGIC_RES[1])
         );
  OAI22_X1 U406 ( .A1(n109), .A2(n189), .B1(n110), .B2(n66), .ZN(LOGIC_RES[2])
         );
  OAI22_X1 U407 ( .A1(n147), .A2(n86), .B1(n148), .B2(n47), .ZN(LOGIC_RES[12])
         );
  OAI22_X1 U408 ( .A1(n139), .A2(n174), .B1(n140), .B2(n51), .ZN(LOGIC_RES[16]) );
  OAI22_X1 U409 ( .A1(n129), .A2(n179), .B1(n130), .B2(n56), .ZN(LOGIC_RES[20]) );
  OAI22_X1 U410 ( .A1(n121), .A2(n183), .B1(n122), .B2(n60), .ZN(LOGIC_RES[24]) );
  OAI22_X1 U411 ( .A1(n113), .A2(n187), .B1(n114), .B2(n64), .ZN(LOGIC_RES[28]) );
  INV_X1 U412 ( .A(OP1[16]), .ZN(n51) );
  INV_X1 U413 ( .A(OP1[17]), .ZN(n52) );
  INV_X1 U414 ( .A(OP1[18]), .ZN(n53) );
  INV_X1 U415 ( .A(OP1[19]), .ZN(n54) );
  INV_X1 U416 ( .A(OP1[20]), .ZN(n56) );
  INV_X1 U417 ( .A(OP1[21]), .ZN(n57) );
  INV_X1 U418 ( .A(OP1[22]), .ZN(n58) );
  INV_X1 U419 ( .A(OP1[23]), .ZN(n59) );
  INV_X1 U420 ( .A(OP1[24]), .ZN(n60) );
  INV_X1 U421 ( .A(OP1[25]), .ZN(n61) );
  INV_X1 U422 ( .A(OP1[26]), .ZN(n62) );
  INV_X1 U423 ( .A(OP1[27]), .ZN(n63) );
  INV_X1 U424 ( .A(OP1[28]), .ZN(n64) );
  INV_X1 U425 ( .A(OP1[29]), .ZN(n65) );
  INV_X1 U426 ( .A(OP1[30]), .ZN(n67) );
  INV_X1 U433 ( .A(OP1[31]), .ZN(n68) );
  NAND2_X1 U437 ( .A1(n157), .A2(n204), .ZN(LOGIC_ARITH) );
  INV_X1 U438 ( .A(LEFT_RIGHT), .ZN(n204) );
  INV_X1 U439 ( .A(n84), .ZN(n205) );
  INV_X1 U440 ( .A(n87), .ZN(n203) );
  INV_X1 U441 ( .A(n80), .ZN(n202) );
  NOR3_X1 U442 ( .A1(n209), .A2(ALU_OPC[3]), .A3(n207), .ZN(n162) );
  NOR3_X1 U443 ( .A1(ALU_OPC[3]), .A2(ALU_OPC[4]), .A3(ALU_OPC[2]), .ZN(n80)
         );
  NAND4_X1 U444 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[1]), .A3(n209), .A4(n206), .ZN(
        n88) );
  NAND4_X1 U445 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[3]), .A3(ALU_OPC[2]), .A4(n201), 
        .ZN(n89) );
  INV_X1 U446 ( .A(ALU_OPC[1]), .ZN(n208) );
  NAND2_X1 U447 ( .A1(n158), .A2(n35), .ZN(LEFT_RIGHT) );
  NOR3_X1 U448 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[4]), .A3(ALU_OPC[2]), .ZN(n156)
         );
  NAND4_X1 U449 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[3]), .A3(n161), .A4(n209), .ZN(
        n157) );
  NOR2_X1 U450 ( .A1(ALU_OPC[4]), .A2(ALU_OPC[2]), .ZN(n161) );
  INV_X1 U451 ( .A(ALU_OPC[2]), .ZN(n207) );
  INV_X1 U452 ( .A(ALU_OPC[3]), .ZN(n206) );
  OAI211_X1 U453 ( .C1(n166), .C2(n167), .A(n206), .B(ALU_OPC[4]), .ZN(n87) );
  NOR2_X1 U454 ( .A1(ALU_OPC[2]), .A2(n208), .ZN(n167) );
  NOR3_X1 U455 ( .A1(n207), .A2(ALU_OPC[1]), .A3(ALU_OPC[0]), .ZN(n166) );
  AND3_X1 U456 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[0]), .A3(n155), .ZN(n92) );
  NOR3_X1 U457 ( .A1(n207), .A2(ALU_OPC[4]), .A3(ALU_OPC[3]), .ZN(n155) );
  INV_X1 U458 ( .A(ALU_OPC[4]), .ZN(n201) );
  INV_X1 U459 ( .A(ALU_OPC[0]), .ZN(n209) );
  OAI21_X1 U460 ( .B1(n78), .B2(n206), .A(n79), .ZN(select_zero_sig) );
  AOI21_X1 U461 ( .B1(ALU_OPC[2]), .B2(n208), .A(ALU_OPC[4]), .ZN(n78) );
  NAND2_X1 U462 ( .A1(n165), .A2(n89), .ZN(OPSel[1]) );
  NAND4_X1 U463 ( .A1(ALU_OPC[4]), .A2(n208), .A3(n207), .A4(n206), .ZN(n165)
         );
  NAND2_X1 U464 ( .A1(n80), .A2(n169), .ZN(n159) );
  XNOR2_X1 U465 ( .A(n208), .B(ALU_OPC[0]), .ZN(n169) );
  AND4_X1 U466 ( .A1(n164), .A2(n88), .A3(n87), .A4(n200), .ZN(n83) );
  INV_X1 U467 ( .A(OPSel[1]), .ZN(n200) );
  OR4_X1 U468 ( .A1(n208), .A2(n207), .A3(ALU_OPC[3]), .A4(ALU_OPC[4]), .ZN(n3) );
  AND2_X1 U469 ( .A1(n160), .A2(n157), .ZN(n81) );
  NAND4_X1 U470 ( .A1(ALU_OPC[0]), .A2(ALU_OPC[3]), .A3(n207), .A4(n201), .ZN(
        n160) );
  NOR3_X1 U471 ( .A1(ALU_OPC[1]), .A2(ALU_OPC[4]), .A3(ALU_OPC[3]), .ZN(n163)
         );
  CLKBUF_X1 U472 ( .A(n205), .Z(n12) );
  CLKBUF_X1 U473 ( .A(n92), .Z(n24) );
  CLKBUF_X1 U474 ( .A(n83), .Z(n34) );
  CLKBUF_X1 U475 ( .A(n81), .Z(n43) );
endmodule


module regn_N32_5 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_4 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N5_2 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 DOUT_reg_4_ ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21) );
  DFFR_X1 DOUT_reg_3_ ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22) );
  DFFR_X1 DOUT_reg_2_ ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23) );
  DFFR_X1 DOUT_reg_1_ ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24) );
  DFFR_X1 DOUT_reg_0_ ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U3 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U4 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U5 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U6 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U7 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U8 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U9 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
  OAI21_X1 U10 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U11 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
endmodule


module regn_N32_3 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module regn_N32_2 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  BUF_X1 U2 ( .A(RST), .Z(n97) );
  BUF_X1 U3 ( .A(RST), .Z(n98) );
  BUF_X1 U4 ( .A(RST), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
endmodule


module Execute_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;
  assign SUM[1] = B[1];
  assign SUM[0] = B[0];

  XNOR2_X1 U1 ( .A(B[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(B[30]), .A2(n56), .ZN(n57) );
  INV_X1 U3 ( .A(B[2]), .ZN(SUM[2]) );
  XOR2_X1 U4 ( .A(B[3]), .B(B[2]), .Z(SUM[3]) );
  XOR2_X1 U5 ( .A(B[4]), .B(n30), .Z(SUM[4]) );
  XOR2_X1 U6 ( .A(B[5]), .B(n31), .Z(SUM[5]) );
  XOR2_X1 U7 ( .A(B[6]), .B(n32), .Z(SUM[6]) );
  XOR2_X1 U8 ( .A(B[7]), .B(n33), .Z(SUM[7]) );
  XOR2_X1 U9 ( .A(B[8]), .B(n34), .Z(SUM[8]) );
  XOR2_X1 U10 ( .A(B[9]), .B(n35), .Z(SUM[9]) );
  XOR2_X1 U11 ( .A(B[10]), .B(n36), .Z(SUM[10]) );
  XOR2_X1 U12 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  XOR2_X1 U13 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  XOR2_X1 U14 ( .A(B[13]), .B(n39), .Z(SUM[13]) );
  XOR2_X1 U15 ( .A(B[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U16 ( .A(B[15]), .B(n41), .Z(SUM[15]) );
  XOR2_X1 U17 ( .A(B[16]), .B(n42), .Z(SUM[16]) );
  XOR2_X1 U18 ( .A(B[17]), .B(n43), .Z(SUM[17]) );
  XOR2_X1 U19 ( .A(B[18]), .B(n44), .Z(SUM[18]) );
  XOR2_X1 U20 ( .A(B[19]), .B(n45), .Z(SUM[19]) );
  XOR2_X1 U21 ( .A(B[20]), .B(n46), .Z(SUM[20]) );
  XOR2_X1 U22 ( .A(B[21]), .B(n47), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(B[22]), .B(n48), .Z(SUM[22]) );
  XOR2_X1 U24 ( .A(B[23]), .B(n49), .Z(SUM[23]) );
  XOR2_X1 U25 ( .A(B[24]), .B(n50), .Z(SUM[24]) );
  XOR2_X1 U26 ( .A(B[25]), .B(n51), .Z(SUM[25]) );
  XOR2_X1 U27 ( .A(B[26]), .B(n52), .Z(SUM[26]) );
  XOR2_X1 U28 ( .A(B[27]), .B(n53), .Z(SUM[27]) );
  XOR2_X1 U29 ( .A(B[28]), .B(n54), .Z(SUM[28]) );
  XOR2_X1 U30 ( .A(B[29]), .B(n55), .Z(SUM[29]) );
  XOR2_X1 U31 ( .A(B[30]), .B(n56), .Z(SUM[30]) );
  AND2_X1 U32 ( .A1(B[3]), .A2(B[2]), .ZN(n30) );
  AND2_X1 U33 ( .A1(B[4]), .A2(n30), .ZN(n31) );
  AND2_X1 U34 ( .A1(B[5]), .A2(n31), .ZN(n32) );
  AND2_X1 U35 ( .A1(B[6]), .A2(n32), .ZN(n33) );
  AND2_X1 U36 ( .A1(B[7]), .A2(n33), .ZN(n34) );
  AND2_X1 U37 ( .A1(B[8]), .A2(n34), .ZN(n35) );
  AND2_X1 U38 ( .A1(B[9]), .A2(n35), .ZN(n36) );
  AND2_X1 U39 ( .A1(B[10]), .A2(n36), .ZN(n37) );
  AND2_X1 U40 ( .A1(B[11]), .A2(n37), .ZN(n38) );
  AND2_X1 U41 ( .A1(B[12]), .A2(n38), .ZN(n39) );
  AND2_X1 U42 ( .A1(B[13]), .A2(n39), .ZN(n40) );
  AND2_X1 U43 ( .A1(B[14]), .A2(n40), .ZN(n41) );
  AND2_X1 U44 ( .A1(B[15]), .A2(n41), .ZN(n42) );
  AND2_X1 U45 ( .A1(B[16]), .A2(n42), .ZN(n43) );
  AND2_X1 U46 ( .A1(B[17]), .A2(n43), .ZN(n44) );
  AND2_X1 U47 ( .A1(B[18]), .A2(n44), .ZN(n45) );
  AND2_X1 U48 ( .A1(B[19]), .A2(n45), .ZN(n46) );
  AND2_X1 U49 ( .A1(B[20]), .A2(n46), .ZN(n47) );
  AND2_X1 U50 ( .A1(B[21]), .A2(n47), .ZN(n48) );
  AND2_X1 U51 ( .A1(B[22]), .A2(n48), .ZN(n49) );
  AND2_X1 U52 ( .A1(B[23]), .A2(n49), .ZN(n50) );
  AND2_X1 U53 ( .A1(B[24]), .A2(n50), .ZN(n51) );
  AND2_X1 U54 ( .A1(B[25]), .A2(n51), .ZN(n52) );
  AND2_X1 U55 ( .A1(B[26]), .A2(n52), .ZN(n53) );
  AND2_X1 U56 ( .A1(B[27]), .A2(n53), .ZN(n54) );
  AND2_X1 U57 ( .A1(B[28]), .A2(n54), .ZN(n55) );
  AND2_X1 U58 ( .A1(B[29]), .A2(n55), .ZN(n56) );
endmodule


module Execute_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:2] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module Execute ( CLK, RST, MUX_A_SEL, MUX_B_SEL, ALU_OPC, ALU_OUTREG_EN, 
        JUMP_TYPE, PC_IN, A_IN, B_IN, IMM_IN, ADD_WR_IN, ADD_RS1_IN, 
        ADD_RS2_IN, ADD_WR_MEM, ADD_WR_WB, RF_WE_MEM, RF_WE_WB, OP_MEM, OP_WB, 
        PC_SEL, ZERO_FLAG, NPC_ABS, NPC_REL, ALU_RES, B_OUT, ADD_WR_OUT );
  input [1:0] MUX_B_SEL;
  input [4:0] ALU_OPC;
  input [1:0] JUMP_TYPE;
  input [31:0] PC_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] ADD_WR_IN;
  input [4:0] ADD_RS1_IN;
  input [4:0] ADD_RS2_IN;
  input [4:0] ADD_WR_MEM;
  input [4:0] ADD_WR_WB;
  input [31:0] OP_MEM;
  input [31:0] OP_WB;
  output [1:0] PC_SEL;
  output [31:0] NPC_ABS;
  output [31:0] NPC_REL;
  output [31:0] ALU_RES;
  output [31:0] B_OUT;
  output [4:0] ADD_WR_OUT;
  input CLK, RST, MUX_A_SEL, ALU_OUTREG_EN, RF_WE_MEM, RF_WE_WB;
  output ZERO_FLAG;
  wire   sig_RST, sig_ZERO_FLAG, N9, N8, N7, N6, N5, N4, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N11, N10, N1, N0, n1;
  wire   [31:0] sig_NPC_ABS;
  wire   [31:0] sig_NPC_REL;
  wire   [1:0] sig_PC_SEL;
  wire   [1:0] FWDA;
  wire   [1:0] FWDB;
  wire   [31:0] OP2_FW;
  wire   [31:0] sig_OP1;
  wire   [31:0] sig_OP2;
  wire   [31:0] sig_ALU_RES;

  Branch_Cond_Unit_NBIT32 Branch_Cond ( .RST(sig_RST), .A(sig_NPC_ABS), 
        .ALU_OPC(ALU_OPC), .JUMP_TYPE(JUMP_TYPE), .PC_SEL(sig_PC_SEL), .ZERO(
        sig_ZERO_FLAG) );
  ff_1 ff0 ( .D(sig_ZERO_FLAG), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(ZERO_FLAG)
         );
  regn_N2 reg0 ( .DIN(sig_PC_SEL), .CLK(CLK), .EN(1'b1), .RST(RST), .DOUT(
        PC_SEL) );
  FWD_Unit FWD ( .RST(sig_RST), .ADD_RS1(ADD_RS1_IN), .ADD_RS2(ADD_RS2_IN), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE_MEM), 
        .RF_WE_WB(RF_WE_WB), .FWDA(FWDA), .FWDB(FWDB) );
  mux41_NBIT32_0 FW1 ( .A(A_IN), .B(OP_WB), .C(OP_MEM), .D(A_IN), .S(FWDA), 
        .Z(sig_NPC_ABS) );
  mux41_NBIT32_4 FW2 ( .A(B_IN), .B(OP_WB), .C(OP_MEM), .D(B_IN), .S(FWDB), 
        .Z(OP2_FW) );
  mux21_NBIT32_4 muxA ( .A(sig_NPC_ABS), .B(PC_IN), .S(MUX_A_SEL), .Z(sig_OP1)
         );
  mux41_NBIT32_3 muxB ( .A(OP2_FW), .B(IMM_IN), .C({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(MUX_B_SEL), .Z(sig_OP2) );
  ALU_NBIT32 alu0 ( .OP1(sig_OP1), .OP2(sig_OP2), .ALU_OPC(ALU_OPC), .ALU_RES(
        sig_ALU_RES) );
  regn_N32_5 alureg ( .DIN(sig_ALU_RES), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(
        RST), .DOUT(ALU_RES) );
  regn_N32_4 B_reg ( .DIN(OP2_FW), .CLK(CLK), .EN(ALU_OUTREG_EN), .RST(RST), 
        .DOUT(B_OUT) );
  regn_N5_2 ADD_WR_reg ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(1'b1), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_3 NPC_ABS_reg ( .DIN(sig_NPC_ABS), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_ABS) );
  regn_N32_2 NPC_REL_reg ( .DIN(sig_NPC_REL), .CLK(CLK), .EN(ALU_OUTREG_EN), 
        .RST(RST), .DOUT(NPC_REL) );
  Execute_DW01_add_1 add_1_root_add_0_root_add_122_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .B(IMM_IN), .CI(1'b0), .SUM({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0})
         );
  Execute_DW01_add_0 add_0_root_add_0_root_add_122_2 ( .A(PC_IN), .B({N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), 
        .CI(1'b0), .SUM(sig_NPC_REL) );
  NOR2_X1 U3 ( .A1(ZERO_FLAG), .A2(n1), .ZN(sig_RST) );
  INV_X1 U4 ( .A(RST), .ZN(n1) );
endmodule


module ff_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFFR_X1 Q_reg ( .D(n3), .CK(CLK), .RN(RST), .Q(Q), .QN(n2) );
  OAI21_X1 U2 ( .B1(n2), .B2(EN), .A(n1), .ZN(n3) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n1) );
endmodule


module regn_N5_1 ( DIN, CLK, EN, RST, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, EN, RST;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 DOUT_reg_4_ ( .D(n16), .CK(CLK), .RN(RST), .Q(DOUT[4]), .QN(n21) );
  DFFR_X1 DOUT_reg_3_ ( .D(n17), .CK(CLK), .RN(RST), .Q(DOUT[3]), .QN(n22) );
  DFFR_X1 DOUT_reg_2_ ( .D(n18), .CK(CLK), .RN(RST), .Q(DOUT[2]), .QN(n23) );
  DFFR_X1 DOUT_reg_1_ ( .D(n19), .CK(CLK), .RN(RST), .Q(DOUT[1]), .QN(n24) );
  DFFR_X1 DOUT_reg_0_ ( .D(n20), .CK(CLK), .RN(RST), .Q(DOUT[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n25), .B2(EN), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(EN), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(EN), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(EN), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(EN), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n26) );
endmodule


module regn_N32_1 ( DIN, CLK, EN, RST, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, EN, RST;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 DOUT_reg_31_ ( .D(n100), .CK(CLK), .RN(n99), .Q(DOUT[31]), .QN(n132)
         );
  DFFR_X1 DOUT_reg_30_ ( .D(n101), .CK(CLK), .RN(n99), .Q(DOUT[30]), .QN(n133)
         );
  DFFR_X1 DOUT_reg_29_ ( .D(n102), .CK(CLK), .RN(n99), .Q(DOUT[29]), .QN(n134)
         );
  DFFR_X1 DOUT_reg_28_ ( .D(n103), .CK(CLK), .RN(n99), .Q(DOUT[28]), .QN(n135)
         );
  DFFR_X1 DOUT_reg_27_ ( .D(n104), .CK(CLK), .RN(n99), .Q(DOUT[27]), .QN(n136)
         );
  DFFR_X1 DOUT_reg_26_ ( .D(n105), .CK(CLK), .RN(n99), .Q(DOUT[26]), .QN(n137)
         );
  DFFR_X1 DOUT_reg_25_ ( .D(n106), .CK(CLK), .RN(n99), .Q(DOUT[25]), .QN(n138)
         );
  DFFR_X1 DOUT_reg_24_ ( .D(n107), .CK(CLK), .RN(n99), .Q(DOUT[24]), .QN(n139)
         );
  DFFR_X1 DOUT_reg_23_ ( .D(n108), .CK(CLK), .RN(n98), .Q(DOUT[23]), .QN(n140)
         );
  DFFR_X1 DOUT_reg_22_ ( .D(n109), .CK(CLK), .RN(n98), .Q(DOUT[22]), .QN(n141)
         );
  DFFR_X1 DOUT_reg_21_ ( .D(n110), .CK(CLK), .RN(n98), .Q(DOUT[21]), .QN(n142)
         );
  DFFR_X1 DOUT_reg_20_ ( .D(n111), .CK(CLK), .RN(n98), .Q(DOUT[20]), .QN(n143)
         );
  DFFR_X1 DOUT_reg_19_ ( .D(n112), .CK(CLK), .RN(n98), .Q(DOUT[19]), .QN(n144)
         );
  DFFR_X1 DOUT_reg_18_ ( .D(n113), .CK(CLK), .RN(n98), .Q(DOUT[18]), .QN(n145)
         );
  DFFR_X1 DOUT_reg_17_ ( .D(n114), .CK(CLK), .RN(n98), .Q(DOUT[17]), .QN(n146)
         );
  DFFR_X1 DOUT_reg_16_ ( .D(n115), .CK(CLK), .RN(n98), .Q(DOUT[16]), .QN(n147)
         );
  DFFR_X1 DOUT_reg_15_ ( .D(n116), .CK(CLK), .RN(n98), .Q(DOUT[15]), .QN(n148)
         );
  DFFR_X1 DOUT_reg_14_ ( .D(n117), .CK(CLK), .RN(n98), .Q(DOUT[14]), .QN(n149)
         );
  DFFR_X1 DOUT_reg_13_ ( .D(n118), .CK(CLK), .RN(n98), .Q(DOUT[13]), .QN(n150)
         );
  DFFR_X1 DOUT_reg_12_ ( .D(n119), .CK(CLK), .RN(n98), .Q(DOUT[12]), .QN(n151)
         );
  DFFR_X1 DOUT_reg_11_ ( .D(n120), .CK(CLK), .RN(n97), .Q(DOUT[11]), .QN(n152)
         );
  DFFR_X1 DOUT_reg_10_ ( .D(n121), .CK(CLK), .RN(n97), .Q(DOUT[10]), .QN(n153)
         );
  DFFR_X1 DOUT_reg_9_ ( .D(n122), .CK(CLK), .RN(n97), .Q(DOUT[9]), .QN(n154)
         );
  DFFR_X1 DOUT_reg_8_ ( .D(n123), .CK(CLK), .RN(n97), .Q(DOUT[8]), .QN(n155)
         );
  DFFR_X1 DOUT_reg_7_ ( .D(n124), .CK(CLK), .RN(n97), .Q(DOUT[7]), .QN(n156)
         );
  DFFR_X1 DOUT_reg_6_ ( .D(n125), .CK(CLK), .RN(n97), .Q(DOUT[6]), .QN(n157)
         );
  DFFR_X1 DOUT_reg_5_ ( .D(n126), .CK(CLK), .RN(n97), .Q(DOUT[5]), .QN(n158)
         );
  DFFR_X1 DOUT_reg_4_ ( .D(n127), .CK(CLK), .RN(n97), .Q(DOUT[4]), .QN(n159)
         );
  DFFR_X1 DOUT_reg_3_ ( .D(n128), .CK(CLK), .RN(n97), .Q(DOUT[3]), .QN(n160)
         );
  DFFR_X1 DOUT_reg_2_ ( .D(n129), .CK(CLK), .RN(n97), .Q(DOUT[2]), .QN(n161)
         );
  DFFR_X1 DOUT_reg_1_ ( .D(n130), .CK(CLK), .RN(n97), .Q(DOUT[1]), .QN(n162)
         );
  DFFR_X1 DOUT_reg_0_ ( .D(n131), .CK(CLK), .RN(n97), .Q(DOUT[0]), .QN(n163)
         );
  OAI21_X1 U2 ( .B1(n163), .B2(EN), .A(n195), .ZN(n131) );
  NAND2_X1 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n195) );
  OAI21_X1 U4 ( .B1(n162), .B2(EN), .A(n194), .ZN(n130) );
  NAND2_X1 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n194) );
  OAI21_X1 U6 ( .B1(n161), .B2(EN), .A(n193), .ZN(n129) );
  NAND2_X1 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n193) );
  OAI21_X1 U8 ( .B1(n160), .B2(EN), .A(n192), .ZN(n128) );
  NAND2_X1 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n192) );
  OAI21_X1 U10 ( .B1(n159), .B2(EN), .A(n191), .ZN(n127) );
  NAND2_X1 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n191) );
  OAI21_X1 U12 ( .B1(n158), .B2(EN), .A(n190), .ZN(n126) );
  NAND2_X1 U13 ( .A1(DIN[5]), .A2(EN), .ZN(n190) );
  OAI21_X1 U14 ( .B1(n157), .B2(EN), .A(n189), .ZN(n125) );
  NAND2_X1 U15 ( .A1(DIN[6]), .A2(EN), .ZN(n189) );
  OAI21_X1 U16 ( .B1(n156), .B2(EN), .A(n188), .ZN(n124) );
  NAND2_X1 U17 ( .A1(DIN[7]), .A2(EN), .ZN(n188) );
  OAI21_X1 U18 ( .B1(n155), .B2(EN), .A(n187), .ZN(n123) );
  NAND2_X1 U19 ( .A1(DIN[8]), .A2(EN), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n154), .B2(EN), .A(n186), .ZN(n122) );
  NAND2_X1 U21 ( .A1(DIN[9]), .A2(EN), .ZN(n186) );
  OAI21_X1 U22 ( .B1(n153), .B2(EN), .A(n185), .ZN(n121) );
  NAND2_X1 U23 ( .A1(DIN[10]), .A2(EN), .ZN(n185) );
  OAI21_X1 U24 ( .B1(n152), .B2(EN), .A(n184), .ZN(n120) );
  NAND2_X1 U25 ( .A1(DIN[11]), .A2(EN), .ZN(n184) );
  OAI21_X1 U26 ( .B1(n151), .B2(EN), .A(n183), .ZN(n119) );
  NAND2_X1 U27 ( .A1(DIN[12]), .A2(EN), .ZN(n183) );
  OAI21_X1 U28 ( .B1(n150), .B2(EN), .A(n182), .ZN(n118) );
  NAND2_X1 U29 ( .A1(DIN[13]), .A2(EN), .ZN(n182) );
  OAI21_X1 U30 ( .B1(n149), .B2(EN), .A(n181), .ZN(n117) );
  NAND2_X1 U31 ( .A1(DIN[14]), .A2(EN), .ZN(n181) );
  OAI21_X1 U32 ( .B1(n148), .B2(EN), .A(n180), .ZN(n116) );
  NAND2_X1 U33 ( .A1(DIN[15]), .A2(EN), .ZN(n180) );
  OAI21_X1 U34 ( .B1(n147), .B2(EN), .A(n179), .ZN(n115) );
  NAND2_X1 U35 ( .A1(DIN[16]), .A2(EN), .ZN(n179) );
  OAI21_X1 U36 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U37 ( .A1(DIN[17]), .A2(EN), .ZN(n178) );
  OAI21_X1 U38 ( .B1(n145), .B2(EN), .A(n177), .ZN(n113) );
  NAND2_X1 U39 ( .A1(DIN[18]), .A2(EN), .ZN(n177) );
  OAI21_X1 U40 ( .B1(n144), .B2(EN), .A(n176), .ZN(n112) );
  NAND2_X1 U41 ( .A1(DIN[19]), .A2(EN), .ZN(n176) );
  OAI21_X1 U42 ( .B1(n143), .B2(EN), .A(n175), .ZN(n111) );
  NAND2_X1 U43 ( .A1(DIN[20]), .A2(EN), .ZN(n175) );
  OAI21_X1 U44 ( .B1(n142), .B2(EN), .A(n174), .ZN(n110) );
  NAND2_X1 U45 ( .A1(DIN[21]), .A2(EN), .ZN(n174) );
  OAI21_X1 U46 ( .B1(n141), .B2(EN), .A(n173), .ZN(n109) );
  NAND2_X1 U47 ( .A1(DIN[22]), .A2(EN), .ZN(n173) );
  OAI21_X1 U48 ( .B1(n140), .B2(EN), .A(n172), .ZN(n108) );
  NAND2_X1 U49 ( .A1(DIN[23]), .A2(EN), .ZN(n172) );
  OAI21_X1 U50 ( .B1(n139), .B2(EN), .A(n171), .ZN(n107) );
  NAND2_X1 U51 ( .A1(DIN[24]), .A2(EN), .ZN(n171) );
  OAI21_X1 U52 ( .B1(n138), .B2(EN), .A(n170), .ZN(n106) );
  NAND2_X1 U53 ( .A1(DIN[25]), .A2(EN), .ZN(n170) );
  OAI21_X1 U54 ( .B1(n137), .B2(EN), .A(n169), .ZN(n105) );
  NAND2_X1 U55 ( .A1(DIN[26]), .A2(EN), .ZN(n169) );
  OAI21_X1 U56 ( .B1(n136), .B2(EN), .A(n168), .ZN(n104) );
  NAND2_X1 U57 ( .A1(DIN[27]), .A2(EN), .ZN(n168) );
  OAI21_X1 U58 ( .B1(n135), .B2(EN), .A(n167), .ZN(n103) );
  NAND2_X1 U59 ( .A1(DIN[28]), .A2(EN), .ZN(n167) );
  OAI21_X1 U60 ( .B1(n134), .B2(EN), .A(n166), .ZN(n102) );
  NAND2_X1 U61 ( .A1(DIN[29]), .A2(EN), .ZN(n166) );
  OAI21_X1 U62 ( .B1(n133), .B2(EN), .A(n165), .ZN(n101) );
  NAND2_X1 U63 ( .A1(DIN[30]), .A2(EN), .ZN(n165) );
  OAI21_X1 U64 ( .B1(n132), .B2(EN), .A(n164), .ZN(n100) );
  NAND2_X1 U65 ( .A1(DIN[31]), .A2(EN), .ZN(n164) );
  BUF_X1 U66 ( .A(RST), .Z(n97) );
  BUF_X1 U67 ( .A(RST), .Z(n98) );
  BUF_X1 U68 ( .A(RST), .Z(n99) );
endmodule


module mux41_NBIT32_2 ( A, B, C, D, S, Z );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Z;
  wire   n1, n4, n5, n6, n7, n20, n21, n22, n23, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n48, n49, n50, n51, n52, n53, n54, n55, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114;

  AND2_X1 U1 ( .A1(S[1]), .A2(n34), .ZN(n1) );
  AND2_X1 U2 ( .A1(S[0]), .A2(n33), .ZN(n4) );
  AND2_X1 U3 ( .A1(n33), .A2(n34), .ZN(n5) );
  AND2_X1 U4 ( .A1(S[0]), .A2(S[1]), .ZN(n6) );
  BUF_X1 U5 ( .A(n5), .Z(n27) );
  BUF_X1 U6 ( .A(n5), .Z(n28) );
  BUF_X1 U7 ( .A(n5), .Z(n29) );
  BUF_X1 U8 ( .A(n1), .Z(n7) );
  BUF_X1 U9 ( .A(n4), .Z(n31) );
  BUF_X1 U10 ( .A(n4), .Z(n30) );
  BUF_X1 U11 ( .A(n1), .Z(n20) );
  BUF_X1 U12 ( .A(n4), .Z(n32) );
  BUF_X1 U13 ( .A(n1), .Z(n21) );
  BUF_X1 U14 ( .A(n6), .Z(n22) );
  BUF_X1 U15 ( .A(n6), .Z(n23) );
  BUF_X1 U16 ( .A(n6), .Z(n26) );
  NAND2_X1 U17 ( .A1(n88), .A2(n87), .ZN(Z[11]) );
  AOI22_X1 U18 ( .A1(D[11]), .A2(n22), .B1(C[11]), .B2(n7), .ZN(n87) );
  AOI22_X1 U19 ( .A1(B[11]), .A2(n30), .B1(A[11]), .B2(n27), .ZN(n88) );
  NAND2_X1 U20 ( .A1(n106), .A2(n105), .ZN(Z[5]) );
  AOI22_X1 U21 ( .A1(D[5]), .A2(n22), .B1(C[5]), .B2(n7), .ZN(n105) );
  AOI22_X1 U22 ( .A1(B[5]), .A2(n30), .B1(A[5]), .B2(n27), .ZN(n106) );
  NAND2_X1 U23 ( .A1(n112), .A2(n111), .ZN(Z[8]) );
  AOI22_X1 U24 ( .A1(D[8]), .A2(n23), .B1(C[8]), .B2(n20), .ZN(n111) );
  AOI22_X1 U25 ( .A1(B[8]), .A2(n31), .B1(A[8]), .B2(n28), .ZN(n112) );
  NAND2_X1 U26 ( .A1(n110), .A2(n109), .ZN(Z[7]) );
  AOI22_X1 U27 ( .A1(D[7]), .A2(n23), .B1(C[7]), .B2(n20), .ZN(n109) );
  AOI22_X1 U28 ( .A1(B[7]), .A2(n31), .B1(A[7]), .B2(n28), .ZN(n110) );
  NAND2_X1 U29 ( .A1(n104), .A2(n103), .ZN(Z[4]) );
  AOI22_X1 U30 ( .A1(D[4]), .A2(n22), .B1(C[4]), .B2(n7), .ZN(n103) );
  AOI22_X1 U31 ( .A1(B[4]), .A2(n30), .B1(A[4]), .B2(n27), .ZN(n104) );
  AOI22_X1 U32 ( .A1(D[15]), .A2(n22), .B1(C[15]), .B2(n7), .ZN(n95) );
  NAND2_X1 U33 ( .A1(n108), .A2(n107), .ZN(Z[6]) );
  AOI22_X1 U34 ( .A1(D[6]), .A2(n23), .B1(C[6]), .B2(n20), .ZN(n107) );
  AOI22_X1 U35 ( .A1(B[6]), .A2(n31), .B1(A[6]), .B2(n28), .ZN(n108) );
  NAND2_X1 U36 ( .A1(n114), .A2(n113), .ZN(Z[9]) );
  AOI22_X1 U37 ( .A1(D[9]), .A2(n23), .B1(C[9]), .B2(n20), .ZN(n113) );
  AOI22_X1 U38 ( .A1(B[9]), .A2(n31), .B1(A[9]), .B2(n28), .ZN(n114) );
  NAND2_X1 U39 ( .A1(n92), .A2(n91), .ZN(Z[13]) );
  AOI22_X1 U40 ( .A1(D[13]), .A2(n22), .B1(C[13]), .B2(n7), .ZN(n91) );
  AOI22_X1 U41 ( .A1(B[13]), .A2(n30), .B1(A[13]), .B2(n27), .ZN(n92) );
  NAND2_X1 U42 ( .A1(n94), .A2(n93), .ZN(Z[14]) );
  AOI22_X1 U43 ( .A1(D[14]), .A2(n22), .B1(C[14]), .B2(n7), .ZN(n93) );
  AOI22_X1 U44 ( .A1(B[14]), .A2(n30), .B1(A[14]), .B2(n27), .ZN(n94) );
  NAND2_X1 U45 ( .A1(n84), .A2(n83), .ZN(Z[0]) );
  AOI22_X1 U46 ( .A1(B[0]), .A2(n30), .B1(A[0]), .B2(n27), .ZN(n84) );
  AOI22_X1 U47 ( .A1(D[0]), .A2(n22), .B1(C[0]), .B2(n7), .ZN(n83) );
  NAND2_X1 U48 ( .A1(n98), .A2(n97), .ZN(Z[1]) );
  AOI22_X1 U49 ( .A1(B[1]), .A2(n30), .B1(A[1]), .B2(n27), .ZN(n98) );
  AOI22_X1 U50 ( .A1(D[1]), .A2(n22), .B1(C[1]), .B2(n7), .ZN(n97) );
  NAND2_X1 U51 ( .A1(n100), .A2(n99), .ZN(Z[2]) );
  AOI22_X1 U52 ( .A1(B[2]), .A2(n30), .B1(A[2]), .B2(n27), .ZN(n100) );
  AOI22_X1 U53 ( .A1(D[2]), .A2(n22), .B1(C[2]), .B2(n7), .ZN(n99) );
  NAND2_X1 U54 ( .A1(n102), .A2(n101), .ZN(Z[3]) );
  AOI22_X1 U55 ( .A1(B[3]), .A2(n30), .B1(A[3]), .B2(n27), .ZN(n102) );
  AOI22_X1 U56 ( .A1(D[3]), .A2(n22), .B1(C[3]), .B2(n7), .ZN(n101) );
  NAND2_X1 U57 ( .A1(n86), .A2(n85), .ZN(Z[10]) );
  AOI22_X1 U58 ( .A1(D[10]), .A2(n22), .B1(C[10]), .B2(n7), .ZN(n85) );
  AOI22_X1 U59 ( .A1(B[10]), .A2(n30), .B1(A[10]), .B2(n27), .ZN(n86) );
  NAND2_X1 U60 ( .A1(n90), .A2(n89), .ZN(Z[12]) );
  AOI22_X1 U61 ( .A1(D[12]), .A2(n22), .B1(C[12]), .B2(n7), .ZN(n89) );
  AOI22_X1 U62 ( .A1(B[12]), .A2(n30), .B1(A[12]), .B2(n27), .ZN(n90) );
  NAND2_X1 U63 ( .A1(n96), .A2(n95), .ZN(Z[15]) );
  AOI22_X1 U64 ( .A1(B[15]), .A2(n30), .B1(A[15]), .B2(n27), .ZN(n96) );
  INV_X1 U65 ( .A(S[1]), .ZN(n33) );
  INV_X1 U66 ( .A(S[0]), .ZN(n34) );
  AOI22_X1 U67 ( .A1(B[16]), .A2(n32), .B1(A[16]), .B2(n29), .ZN(n36) );
  AOI22_X1 U68 ( .A1(D[16]), .A2(n26), .B1(C[16]), .B2(n21), .ZN(n35) );
  NAND2_X1 U69 ( .A1(n36), .A2(n35), .ZN(Z[16]) );
  AOI22_X1 U70 ( .A1(B[17]), .A2(n32), .B1(A[17]), .B2(n29), .ZN(n38) );
  AOI22_X1 U71 ( .A1(D[17]), .A2(n26), .B1(C[17]), .B2(n21), .ZN(n37) );
  NAND2_X1 U72 ( .A1(n38), .A2(n37), .ZN(Z[17]) );
  AOI22_X1 U73 ( .A1(B[18]), .A2(n32), .B1(A[18]), .B2(n29), .ZN(n40) );
  AOI22_X1 U74 ( .A1(D[18]), .A2(n26), .B1(C[18]), .B2(n21), .ZN(n39) );
  NAND2_X1 U75 ( .A1(n40), .A2(n39), .ZN(Z[18]) );
  AOI22_X1 U76 ( .A1(B[19]), .A2(n31), .B1(A[19]), .B2(n28), .ZN(n42) );
  AOI22_X1 U77 ( .A1(D[19]), .A2(n23), .B1(C[19]), .B2(n20), .ZN(n41) );
  NAND2_X1 U78 ( .A1(n42), .A2(n41), .ZN(Z[19]) );
  AOI22_X1 U79 ( .A1(B[20]), .A2(n31), .B1(A[20]), .B2(n28), .ZN(n44) );
  AOI22_X1 U80 ( .A1(D[20]), .A2(n23), .B1(C[20]), .B2(n20), .ZN(n43) );
  NAND2_X1 U81 ( .A1(n44), .A2(n43), .ZN(Z[20]) );
  AOI22_X1 U82 ( .A1(B[21]), .A2(n31), .B1(A[21]), .B2(n28), .ZN(n48) );
  AOI22_X1 U83 ( .A1(D[21]), .A2(n23), .B1(C[21]), .B2(n20), .ZN(n45) );
  NAND2_X1 U84 ( .A1(n48), .A2(n45), .ZN(Z[21]) );
  AOI22_X1 U85 ( .A1(B[22]), .A2(n31), .B1(A[22]), .B2(n28), .ZN(n50) );
  AOI22_X1 U86 ( .A1(D[22]), .A2(n23), .B1(C[22]), .B2(n20), .ZN(n49) );
  NAND2_X1 U87 ( .A1(n50), .A2(n49), .ZN(Z[22]) );
  AOI22_X1 U88 ( .A1(B[23]), .A2(n31), .B1(A[23]), .B2(n28), .ZN(n52) );
  AOI22_X1 U89 ( .A1(D[23]), .A2(n23), .B1(C[23]), .B2(n20), .ZN(n51) );
  NAND2_X1 U90 ( .A1(n52), .A2(n51), .ZN(Z[23]) );
  AOI22_X1 U91 ( .A1(B[24]), .A2(n31), .B1(A[24]), .B2(n28), .ZN(n54) );
  AOI22_X1 U92 ( .A1(D[24]), .A2(n23), .B1(C[24]), .B2(n20), .ZN(n53) );
  NAND2_X1 U93 ( .A1(n54), .A2(n53), .ZN(Z[24]) );
  AOI22_X1 U94 ( .A1(B[25]), .A2(n31), .B1(A[25]), .B2(n28), .ZN(n70) );
  AOI22_X1 U95 ( .A1(D[25]), .A2(n23), .B1(C[25]), .B2(n20), .ZN(n55) );
  NAND2_X1 U96 ( .A1(n70), .A2(n55), .ZN(Z[25]) );
  AOI22_X1 U97 ( .A1(B[26]), .A2(n31), .B1(A[26]), .B2(n28), .ZN(n72) );
  AOI22_X1 U98 ( .A1(D[26]), .A2(n23), .B1(C[26]), .B2(n20), .ZN(n71) );
  NAND2_X1 U99 ( .A1(n72), .A2(n71), .ZN(Z[26]) );
  AOI22_X1 U100 ( .A1(B[27]), .A2(n31), .B1(A[27]), .B2(n28), .ZN(n74) );
  AOI22_X1 U101 ( .A1(D[27]), .A2(n23), .B1(C[27]), .B2(n20), .ZN(n73) );
  NAND2_X1 U102 ( .A1(n74), .A2(n73), .ZN(Z[27]) );
  AOI22_X1 U103 ( .A1(B[28]), .A2(n31), .B1(A[28]), .B2(n28), .ZN(n76) );
  AOI22_X1 U104 ( .A1(D[28]), .A2(n23), .B1(C[28]), .B2(n20), .ZN(n75) );
  NAND2_X1 U105 ( .A1(n76), .A2(n75), .ZN(Z[28]) );
  AOI22_X1 U106 ( .A1(B[29]), .A2(n31), .B1(A[29]), .B2(n28), .ZN(n78) );
  AOI22_X1 U107 ( .A1(D[29]), .A2(n23), .B1(C[29]), .B2(n20), .ZN(n77) );
  NAND2_X1 U108 ( .A1(n78), .A2(n77), .ZN(Z[29]) );
  AOI22_X1 U109 ( .A1(B[30]), .A2(n31), .B1(A[30]), .B2(n28), .ZN(n80) );
  AOI22_X1 U110 ( .A1(D[30]), .A2(n23), .B1(C[30]), .B2(n20), .ZN(n79) );
  NAND2_X1 U111 ( .A1(n80), .A2(n79), .ZN(Z[30]) );
  AOI22_X1 U112 ( .A1(B[31]), .A2(n31), .B1(A[31]), .B2(n28), .ZN(n82) );
  AOI22_X1 U113 ( .A1(D[31]), .A2(n23), .B1(C[31]), .B2(n20), .ZN(n81) );
  NAND2_X1 U114 ( .A1(n82), .A2(n81), .ZN(Z[31]) );
endmodule


module Memory ( CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, PC_SEL, NPC_IN, 
        NPC_ABS, NPC_REL, ALU_RES_IN, B_IN, ADD_WR_IN, DRAM_DATA_IN, 
        LOAD_TYPE_IN, STORE_TYPE_IN, PC_OUT, DRAM_R_OUT, DRAM_W_OUT, 
        DRAM_ADDR_OUT, DRAM_DATA_OUT, DATA_OUT, ALU_RES_OUT, OP_MEM, 
        ADD_WR_MEM, ADD_WR_OUT, LOAD_TYPE_OUT, STORE_TYPE_OUT );
  input [1:0] PC_SEL;
  input [31:0] NPC_IN;
  input [31:0] NPC_ABS;
  input [31:0] NPC_REL;
  input [31:0] ALU_RES_IN;
  input [31:0] B_IN;
  input [4:0] ADD_WR_IN;
  input [31:0] DRAM_DATA_IN;
  input [1:0] LOAD_TYPE_IN;
  output [31:0] PC_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DRAM_DATA_OUT;
  output [31:0] DATA_OUT;
  output [31:0] ALU_RES_OUT;
  output [31:0] OP_MEM;
  output [4:0] ADD_WR_MEM;
  output [4:0] ADD_WR_OUT;
  output [1:0] LOAD_TYPE_OUT;
  input CLK, RST, MEM_EN_IN, DRAM_R_IN, DRAM_W_IN, STORE_TYPE_IN;
  output DRAM_R_OUT, DRAM_W_OUT, STORE_TYPE_OUT;
  wire   DRAM_R_IN, DRAM_W_IN, STORE_TYPE_IN;
  assign DRAM_R_OUT = DRAM_R_IN;
  assign DRAM_W_OUT = DRAM_W_IN;
  assign OP_MEM[31] = ALU_RES_IN[31];
  assign DRAM_ADDR_OUT[31] = ALU_RES_IN[31];
  assign OP_MEM[30] = ALU_RES_IN[30];
  assign DRAM_ADDR_OUT[30] = ALU_RES_IN[30];
  assign OP_MEM[29] = ALU_RES_IN[29];
  assign DRAM_ADDR_OUT[29] = ALU_RES_IN[29];
  assign OP_MEM[28] = ALU_RES_IN[28];
  assign DRAM_ADDR_OUT[28] = ALU_RES_IN[28];
  assign OP_MEM[27] = ALU_RES_IN[27];
  assign DRAM_ADDR_OUT[27] = ALU_RES_IN[27];
  assign OP_MEM[26] = ALU_RES_IN[26];
  assign DRAM_ADDR_OUT[26] = ALU_RES_IN[26];
  assign OP_MEM[25] = ALU_RES_IN[25];
  assign DRAM_ADDR_OUT[25] = ALU_RES_IN[25];
  assign OP_MEM[24] = ALU_RES_IN[24];
  assign DRAM_ADDR_OUT[24] = ALU_RES_IN[24];
  assign OP_MEM[23] = ALU_RES_IN[23];
  assign DRAM_ADDR_OUT[23] = ALU_RES_IN[23];
  assign OP_MEM[22] = ALU_RES_IN[22];
  assign DRAM_ADDR_OUT[22] = ALU_RES_IN[22];
  assign OP_MEM[21] = ALU_RES_IN[21];
  assign DRAM_ADDR_OUT[21] = ALU_RES_IN[21];
  assign OP_MEM[20] = ALU_RES_IN[20];
  assign DRAM_ADDR_OUT[20] = ALU_RES_IN[20];
  assign OP_MEM[19] = ALU_RES_IN[19];
  assign DRAM_ADDR_OUT[19] = ALU_RES_IN[19];
  assign OP_MEM[18] = ALU_RES_IN[18];
  assign DRAM_ADDR_OUT[18] = ALU_RES_IN[18];
  assign OP_MEM[17] = ALU_RES_IN[17];
  assign DRAM_ADDR_OUT[17] = ALU_RES_IN[17];
  assign OP_MEM[16] = ALU_RES_IN[16];
  assign DRAM_ADDR_OUT[16] = ALU_RES_IN[16];
  assign OP_MEM[15] = ALU_RES_IN[15];
  assign DRAM_ADDR_OUT[15] = ALU_RES_IN[15];
  assign OP_MEM[14] = ALU_RES_IN[14];
  assign DRAM_ADDR_OUT[14] = ALU_RES_IN[14];
  assign OP_MEM[13] = ALU_RES_IN[13];
  assign DRAM_ADDR_OUT[13] = ALU_RES_IN[13];
  assign OP_MEM[12] = ALU_RES_IN[12];
  assign DRAM_ADDR_OUT[12] = ALU_RES_IN[12];
  assign OP_MEM[11] = ALU_RES_IN[11];
  assign DRAM_ADDR_OUT[11] = ALU_RES_IN[11];
  assign OP_MEM[10] = ALU_RES_IN[10];
  assign DRAM_ADDR_OUT[10] = ALU_RES_IN[10];
  assign OP_MEM[9] = ALU_RES_IN[9];
  assign DRAM_ADDR_OUT[9] = ALU_RES_IN[9];
  assign OP_MEM[8] = ALU_RES_IN[8];
  assign DRAM_ADDR_OUT[8] = ALU_RES_IN[8];
  assign OP_MEM[7] = ALU_RES_IN[7];
  assign DRAM_ADDR_OUT[7] = ALU_RES_IN[7];
  assign OP_MEM[6] = ALU_RES_IN[6];
  assign DRAM_ADDR_OUT[6] = ALU_RES_IN[6];
  assign OP_MEM[5] = ALU_RES_IN[5];
  assign DRAM_ADDR_OUT[5] = ALU_RES_IN[5];
  assign OP_MEM[4] = ALU_RES_IN[4];
  assign DRAM_ADDR_OUT[4] = ALU_RES_IN[4];
  assign OP_MEM[3] = ALU_RES_IN[3];
  assign DRAM_ADDR_OUT[3] = ALU_RES_IN[3];
  assign OP_MEM[2] = ALU_RES_IN[2];
  assign DRAM_ADDR_OUT[2] = ALU_RES_IN[2];
  assign OP_MEM[1] = ALU_RES_IN[1];
  assign DRAM_ADDR_OUT[1] = ALU_RES_IN[1];
  assign OP_MEM[0] = ALU_RES_IN[0];
  assign DRAM_ADDR_OUT[0] = ALU_RES_IN[0];
  assign DRAM_DATA_OUT[31] = B_IN[31];
  assign DRAM_DATA_OUT[30] = B_IN[30];
  assign DRAM_DATA_OUT[29] = B_IN[29];
  assign DRAM_DATA_OUT[28] = B_IN[28];
  assign DRAM_DATA_OUT[27] = B_IN[27];
  assign DRAM_DATA_OUT[26] = B_IN[26];
  assign DRAM_DATA_OUT[25] = B_IN[25];
  assign DRAM_DATA_OUT[24] = B_IN[24];
  assign DRAM_DATA_OUT[23] = B_IN[23];
  assign DRAM_DATA_OUT[22] = B_IN[22];
  assign DRAM_DATA_OUT[21] = B_IN[21];
  assign DRAM_DATA_OUT[20] = B_IN[20];
  assign DRAM_DATA_OUT[19] = B_IN[19];
  assign DRAM_DATA_OUT[18] = B_IN[18];
  assign DRAM_DATA_OUT[17] = B_IN[17];
  assign DRAM_DATA_OUT[16] = B_IN[16];
  assign DRAM_DATA_OUT[15] = B_IN[15];
  assign DRAM_DATA_OUT[14] = B_IN[14];
  assign DRAM_DATA_OUT[13] = B_IN[13];
  assign DRAM_DATA_OUT[12] = B_IN[12];
  assign DRAM_DATA_OUT[11] = B_IN[11];
  assign DRAM_DATA_OUT[10] = B_IN[10];
  assign DRAM_DATA_OUT[9] = B_IN[9];
  assign DRAM_DATA_OUT[8] = B_IN[8];
  assign DRAM_DATA_OUT[7] = B_IN[7];
  assign DRAM_DATA_OUT[6] = B_IN[6];
  assign DRAM_DATA_OUT[5] = B_IN[5];
  assign DRAM_DATA_OUT[4] = B_IN[4];
  assign DRAM_DATA_OUT[3] = B_IN[3];
  assign DRAM_DATA_OUT[2] = B_IN[2];
  assign DRAM_DATA_OUT[1] = B_IN[1];
  assign DRAM_DATA_OUT[0] = B_IN[0];
  assign DATA_OUT[31] = DRAM_DATA_IN[31];
  assign DATA_OUT[30] = DRAM_DATA_IN[30];
  assign DATA_OUT[29] = DRAM_DATA_IN[29];
  assign DATA_OUT[28] = DRAM_DATA_IN[28];
  assign DATA_OUT[27] = DRAM_DATA_IN[27];
  assign DATA_OUT[26] = DRAM_DATA_IN[26];
  assign DATA_OUT[25] = DRAM_DATA_IN[25];
  assign DATA_OUT[24] = DRAM_DATA_IN[24];
  assign DATA_OUT[23] = DRAM_DATA_IN[23];
  assign DATA_OUT[22] = DRAM_DATA_IN[22];
  assign DATA_OUT[21] = DRAM_DATA_IN[21];
  assign DATA_OUT[20] = DRAM_DATA_IN[20];
  assign DATA_OUT[19] = DRAM_DATA_IN[19];
  assign DATA_OUT[18] = DRAM_DATA_IN[18];
  assign DATA_OUT[17] = DRAM_DATA_IN[17];
  assign DATA_OUT[16] = DRAM_DATA_IN[16];
  assign DATA_OUT[15] = DRAM_DATA_IN[15];
  assign DATA_OUT[14] = DRAM_DATA_IN[14];
  assign DATA_OUT[13] = DRAM_DATA_IN[13];
  assign DATA_OUT[12] = DRAM_DATA_IN[12];
  assign DATA_OUT[11] = DRAM_DATA_IN[11];
  assign DATA_OUT[10] = DRAM_DATA_IN[10];
  assign DATA_OUT[9] = DRAM_DATA_IN[9];
  assign DATA_OUT[8] = DRAM_DATA_IN[8];
  assign DATA_OUT[7] = DRAM_DATA_IN[7];
  assign DATA_OUT[6] = DRAM_DATA_IN[6];
  assign DATA_OUT[5] = DRAM_DATA_IN[5];
  assign DATA_OUT[4] = DRAM_DATA_IN[4];
  assign DATA_OUT[3] = DRAM_DATA_IN[3];
  assign DATA_OUT[2] = DRAM_DATA_IN[2];
  assign DATA_OUT[1] = DRAM_DATA_IN[1];
  assign DATA_OUT[0] = DRAM_DATA_IN[0];
  assign ADD_WR_MEM[4] = ADD_WR_IN[4];
  assign ADD_WR_MEM[3] = ADD_WR_IN[3];
  assign ADD_WR_MEM[2] = ADD_WR_IN[2];
  assign ADD_WR_MEM[1] = ADD_WR_IN[1];
  assign ADD_WR_MEM[0] = ADD_WR_IN[0];
  assign LOAD_TYPE_OUT[1] = LOAD_TYPE_IN[1];
  assign LOAD_TYPE_OUT[0] = LOAD_TYPE_IN[0];
  assign STORE_TYPE_OUT = STORE_TYPE_IN;

  regn_N5_1 reg0 ( .DIN(ADD_WR_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ADD_WR_OUT) );
  regn_N32_1 reg1 ( .DIN(ALU_RES_IN), .CLK(CLK), .EN(MEM_EN_IN), .RST(RST), 
        .DOUT(ALU_RES_OUT) );
  mux41_NBIT32_2 PCsel ( .A(NPC_IN), .B(NPC_REL), .C(NPC_ABS), .D({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(PC_SEL), .Z(PC_OUT) );
endmodule


module ff_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n4, n5, n6;

  DFFR_X1 Q_reg ( .D(n4), .CK(CLK), .RN(RST), .Q(Q), .QN(n5) );
  OAI21_X1 U2 ( .B1(n5), .B2(EN), .A(n6), .ZN(n4) );
  NAND2_X1 U3 ( .A1(EN), .A2(D), .ZN(n6) );
endmodule


module mux21_NBIT32_3 ( A, B, S, Z );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Z;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n80), .ZN(Z[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n1), .B1(B[1]), .B2(S), .ZN(n80) );
  INV_X1 U6 ( .A(n69), .ZN(Z[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(S), .ZN(n69) );
  INV_X1 U8 ( .A(n94), .ZN(Z[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n3), .B1(B[3]), .B2(S), .ZN(n94) );
  INV_X1 U10 ( .A(n81), .ZN(Z[20]) );
  AOI22_X1 U11 ( .A1(A[20]), .A2(n2), .B1(B[20]), .B2(S), .ZN(n81) );
  INV_X1 U12 ( .A(n82), .ZN(Z[21]) );
  AOI22_X1 U13 ( .A1(A[21]), .A2(n2), .B1(B[21]), .B2(S), .ZN(n82) );
  INV_X1 U14 ( .A(n83), .ZN(Z[22]) );
  AOI22_X1 U15 ( .A1(A[22]), .A2(n2), .B1(B[22]), .B2(S), .ZN(n83) );
  INV_X1 U16 ( .A(n84), .ZN(Z[23]) );
  AOI22_X1 U17 ( .A1(A[23]), .A2(n2), .B1(B[23]), .B2(S), .ZN(n84) );
  INV_X1 U18 ( .A(n77), .ZN(Z[17]) );
  AOI22_X1 U19 ( .A1(A[17]), .A2(n1), .B1(B[17]), .B2(S), .ZN(n77) );
  INV_X1 U20 ( .A(n78), .ZN(Z[18]) );
  AOI22_X1 U21 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(S), .ZN(n78) );
  INV_X1 U22 ( .A(n79), .ZN(Z[19]) );
  AOI22_X1 U23 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(S), .ZN(n79) );
  INV_X1 U24 ( .A(n73), .ZN(Z[13]) );
  AOI22_X1 U25 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(S), .ZN(n73) );
  INV_X1 U26 ( .A(n74), .ZN(Z[14]) );
  AOI22_X1 U27 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(S), .ZN(n74) );
  INV_X1 U28 ( .A(n75), .ZN(Z[15]) );
  AOI22_X1 U29 ( .A1(A[15]), .A2(n1), .B1(B[15]), .B2(S), .ZN(n75) );
  INV_X1 U30 ( .A(n76), .ZN(Z[16]) );
  AOI22_X1 U31 ( .A1(A[16]), .A2(n1), .B1(B[16]), .B2(S), .ZN(n76) );
  INV_X1 U32 ( .A(n70), .ZN(Z[10]) );
  AOI22_X1 U33 ( .A1(A[10]), .A2(n1), .B1(B[10]), .B2(S), .ZN(n70) );
  INV_X1 U34 ( .A(n71), .ZN(Z[11]) );
  AOI22_X1 U35 ( .A1(A[11]), .A2(n1), .B1(B[11]), .B2(S), .ZN(n71) );
  INV_X1 U36 ( .A(n72), .ZN(Z[12]) );
  AOI22_X1 U37 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(S), .ZN(n72) );
  INV_X1 U38 ( .A(n97), .ZN(Z[6]) );
  AOI22_X1 U39 ( .A1(A[6]), .A2(n3), .B1(B[6]), .B2(S), .ZN(n97) );
  INV_X1 U40 ( .A(n98), .ZN(Z[7]) );
  AOI22_X1 U41 ( .A1(A[7]), .A2(n3), .B1(B[7]), .B2(S), .ZN(n98) );
  INV_X1 U42 ( .A(n99), .ZN(Z[8]) );
  AOI22_X1 U43 ( .A1(A[8]), .A2(n3), .B1(B[8]), .B2(S), .ZN(n99) );
  INV_X1 U44 ( .A(n95), .ZN(Z[4]) );
  AOI22_X1 U45 ( .A1(A[4]), .A2(n3), .B1(B[4]), .B2(S), .ZN(n95) );
  INV_X1 U46 ( .A(n96), .ZN(Z[5]) );
  AOI22_X1 U47 ( .A1(A[5]), .A2(n3), .B1(B[5]), .B2(S), .ZN(n96) );
  INV_X1 U48 ( .A(n89), .ZN(Z[28]) );
  AOI22_X1 U49 ( .A1(A[28]), .A2(n2), .B1(B[28]), .B2(S), .ZN(n89) );
  INV_X1 U50 ( .A(n90), .ZN(Z[29]) );
  AOI22_X1 U51 ( .A1(A[29]), .A2(n2), .B1(B[29]), .B2(S), .ZN(n90) );
  INV_X1 U52 ( .A(n91), .ZN(Z[2]) );
  AOI22_X1 U53 ( .A1(A[2]), .A2(n2), .B1(B[2]), .B2(S), .ZN(n91) );
  INV_X1 U54 ( .A(n92), .ZN(Z[30]) );
  AOI22_X1 U55 ( .A1(A[30]), .A2(n2), .B1(B[30]), .B2(S), .ZN(n92) );
  INV_X1 U56 ( .A(n85), .ZN(Z[24]) );
  AOI22_X1 U57 ( .A1(A[24]), .A2(n2), .B1(B[24]), .B2(S), .ZN(n85) );
  INV_X1 U58 ( .A(n86), .ZN(Z[25]) );
  AOI22_X1 U59 ( .A1(A[25]), .A2(n2), .B1(B[25]), .B2(S), .ZN(n86) );
  INV_X1 U60 ( .A(n87), .ZN(Z[26]) );
  AOI22_X1 U61 ( .A1(A[26]), .A2(n2), .B1(B[26]), .B2(S), .ZN(n87) );
  INV_X1 U62 ( .A(n88), .ZN(Z[27]) );
  AOI22_X1 U63 ( .A1(A[27]), .A2(n2), .B1(B[27]), .B2(S), .ZN(n88) );
  INV_X1 U64 ( .A(n93), .ZN(Z[31]) );
  AOI22_X1 U65 ( .A1(A[31]), .A2(n3), .B1(B[31]), .B2(S), .ZN(n93) );
  INV_X1 U66 ( .A(n100), .ZN(Z[9]) );
  AOI22_X1 U67 ( .A1(A[9]), .A2(n3), .B1(S), .B2(B[9]), .ZN(n100) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module Writeback ( WB_MUX_SEL, DATA_IN, ALU_RES_IN, ADD_WR_IN, DATA_OUT, 
        ADD_WR_OUT );
  input [31:0] DATA_IN;
  input [31:0] ALU_RES_IN;
  input [4:0] ADD_WR_IN;
  output [31:0] DATA_OUT;
  output [4:0] ADD_WR_OUT;
  input WB_MUX_SEL;

  assign ADD_WR_OUT[4] = ADD_WR_IN[4];
  assign ADD_WR_OUT[3] = ADD_WR_IN[3];
  assign ADD_WR_OUT[2] = ADD_WR_IN[2];
  assign ADD_WR_OUT[1] = ADD_WR_IN[1];
  assign ADD_WR_OUT[0] = ADD_WR_IN[0];

  mux21_NBIT32_3 WBmux ( .A(ALU_RES_IN), .B(DATA_IN), .S(WB_MUX_SEL), .Z(
        DATA_OUT) );
endmodule


module HazardDetection_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XNOR2_X1 U1 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  XOR2_X1 U2 ( .A(A[30]), .B(n35), .Z(SUM[30]) );
  XOR2_X1 U3 ( .A(A[16]), .B(n21), .Z(SUM[16]) );
  XOR2_X1 U4 ( .A(A[17]), .B(n22), .Z(SUM[17]) );
  XOR2_X1 U5 ( .A(A[18]), .B(n23), .Z(SUM[18]) );
  XOR2_X1 U6 ( .A(A[19]), .B(n24), .Z(SUM[19]) );
  XOR2_X1 U7 ( .A(A[20]), .B(n25), .Z(SUM[20]) );
  XOR2_X1 U8 ( .A(A[21]), .B(n26), .Z(SUM[21]) );
  XOR2_X1 U9 ( .A(A[22]), .B(n27), .Z(SUM[22]) );
  XOR2_X1 U10 ( .A(A[23]), .B(n28), .Z(SUM[23]) );
  XOR2_X1 U11 ( .A(A[24]), .B(n29), .Z(SUM[24]) );
  XOR2_X1 U12 ( .A(A[25]), .B(n30), .Z(SUM[25]) );
  XOR2_X1 U13 ( .A(A[26]), .B(n31), .Z(SUM[26]) );
  XOR2_X1 U14 ( .A(A[27]), .B(n32), .Z(SUM[27]) );
  XOR2_X1 U15 ( .A(A[28]), .B(n33), .Z(SUM[28]) );
  XOR2_X1 U16 ( .A(A[29]), .B(n34), .Z(SUM[29]) );
  NAND2_X1 U17 ( .A1(A[30]), .A2(n35), .ZN(n57) );
  AND2_X1 U18 ( .A1(A[11]), .A2(n43), .ZN(n17) );
  AND2_X1 U19 ( .A1(A[12]), .A2(n17), .ZN(n18) );
  AND2_X1 U20 ( .A1(A[13]), .A2(n18), .ZN(n19) );
  AND2_X1 U21 ( .A1(A[14]), .A2(n19), .ZN(n20) );
  AND2_X1 U22 ( .A1(A[15]), .A2(n20), .ZN(n21) );
  AND2_X1 U23 ( .A1(A[16]), .A2(n21), .ZN(n22) );
  AND2_X1 U24 ( .A1(A[17]), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(A[18]), .A2(n23), .ZN(n24) );
  AND2_X1 U26 ( .A1(A[19]), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[20]), .A2(n25), .ZN(n26) );
  AND2_X1 U28 ( .A1(A[21]), .A2(n26), .ZN(n27) );
  AND2_X1 U29 ( .A1(A[22]), .A2(n27), .ZN(n28) );
  AND2_X1 U30 ( .A1(A[23]), .A2(n28), .ZN(n29) );
  AND2_X1 U31 ( .A1(A[24]), .A2(n29), .ZN(n30) );
  AND2_X1 U32 ( .A1(A[25]), .A2(n30), .ZN(n31) );
  AND2_X1 U33 ( .A1(A[26]), .A2(n31), .ZN(n32) );
  AND2_X1 U34 ( .A1(A[27]), .A2(n32), .ZN(n33) );
  AND2_X1 U35 ( .A1(A[28]), .A2(n33), .ZN(n34) );
  AND2_X1 U36 ( .A1(A[29]), .A2(n34), .ZN(n35) );
  AND2_X1 U37 ( .A1(A[9]), .A2(n42), .ZN(n36) );
  AND2_X1 U38 ( .A1(A[3]), .A2(A[2]), .ZN(n37) );
  AND2_X1 U39 ( .A1(A[4]), .A2(n37), .ZN(n38) );
  AND2_X1 U40 ( .A1(A[5]), .A2(n38), .ZN(n39) );
  AND2_X1 U41 ( .A1(A[6]), .A2(n39), .ZN(n40) );
  AND2_X1 U42 ( .A1(A[7]), .A2(n40), .ZN(n41) );
  AND2_X1 U43 ( .A1(A[8]), .A2(n41), .ZN(n42) );
  AND2_X1 U44 ( .A1(A[10]), .A2(n36), .ZN(n43) );
  INV_X1 U45 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U46 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U47 ( .A(A[9]), .B(n42), .Z(SUM[9]) );
  XOR2_X1 U48 ( .A(A[11]), .B(n43), .Z(SUM[11]) );
  XOR2_X1 U49 ( .A(A[12]), .B(n17), .Z(SUM[12]) );
  XOR2_X1 U50 ( .A(A[13]), .B(n18), .Z(SUM[13]) );
  XOR2_X1 U51 ( .A(A[14]), .B(n19), .Z(SUM[14]) );
  XOR2_X1 U52 ( .A(A[15]), .B(n20), .Z(SUM[15]) );
  XOR2_X1 U53 ( .A(A[4]), .B(n37), .Z(SUM[4]) );
  XOR2_X1 U54 ( .A(A[5]), .B(n38), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[6]), .B(n39), .Z(SUM[6]) );
  XOR2_X1 U56 ( .A(A[7]), .B(n40), .Z(SUM[7]) );
  XOR2_X1 U57 ( .A(A[8]), .B(n41), .Z(SUM[8]) );
  XOR2_X1 U58 ( .A(A[10]), .B(n36), .Z(SUM[10]) );
endmodule


module HazardDetection ( RST, ADD_RS1, ADD_RS2, ADD_WR, DRAM_R, INS_IN, PC_IN, 
        Bubble, HDU_INS_OUT, HDU_PC_OUT, HDU_NPC_OUT );
  input [4:0] ADD_RS1;
  input [4:0] ADD_RS2;
  input [4:0] ADD_WR;
  input [31:0] INS_IN;
  input [31:0] PC_IN;
  output [31:0] HDU_INS_OUT;
  output [31:0] HDU_PC_OUT;
  output [31:0] HDU_NPC_OUT;
  input RST, DRAM_R;
  output Bubble;
  wire   n1, n2, n3, n4, n5, n6, n9, n10, n12, n13, n14, n15, n16;
  assign HDU_INS_OUT[31] = INS_IN[31];
  assign HDU_INS_OUT[30] = INS_IN[30];
  assign HDU_INS_OUT[29] = INS_IN[29];
  assign HDU_INS_OUT[28] = INS_IN[28];
  assign HDU_INS_OUT[27] = INS_IN[27];
  assign HDU_INS_OUT[26] = INS_IN[26];
  assign HDU_INS_OUT[25] = INS_IN[25];
  assign HDU_INS_OUT[24] = INS_IN[24];
  assign HDU_INS_OUT[23] = INS_IN[23];
  assign HDU_INS_OUT[22] = INS_IN[22];
  assign HDU_INS_OUT[21] = INS_IN[21];
  assign HDU_INS_OUT[20] = INS_IN[20];
  assign HDU_INS_OUT[19] = INS_IN[19];
  assign HDU_INS_OUT[18] = INS_IN[18];
  assign HDU_INS_OUT[17] = INS_IN[17];
  assign HDU_INS_OUT[16] = INS_IN[16];
  assign HDU_INS_OUT[15] = INS_IN[15];
  assign HDU_INS_OUT[14] = INS_IN[14];
  assign HDU_INS_OUT[13] = INS_IN[13];
  assign HDU_INS_OUT[12] = INS_IN[12];
  assign HDU_INS_OUT[11] = INS_IN[11];
  assign HDU_INS_OUT[10] = INS_IN[10];
  assign HDU_INS_OUT[9] = INS_IN[9];
  assign HDU_INS_OUT[8] = INS_IN[8];
  assign HDU_INS_OUT[7] = INS_IN[7];
  assign HDU_INS_OUT[6] = INS_IN[6];
  assign HDU_INS_OUT[5] = INS_IN[5];
  assign HDU_INS_OUT[4] = INS_IN[4];
  assign HDU_INS_OUT[3] = INS_IN[3];
  assign HDU_INS_OUT[2] = INS_IN[2];
  assign HDU_INS_OUT[1] = INS_IN[1];
  assign HDU_INS_OUT[0] = INS_IN[0];
  assign HDU_PC_OUT[31] = PC_IN[31];
  assign HDU_PC_OUT[30] = PC_IN[30];
  assign HDU_PC_OUT[29] = PC_IN[29];
  assign HDU_PC_OUT[28] = PC_IN[28];
  assign HDU_PC_OUT[27] = PC_IN[27];
  assign HDU_PC_OUT[26] = PC_IN[26];
  assign HDU_PC_OUT[25] = PC_IN[25];
  assign HDU_PC_OUT[24] = PC_IN[24];
  assign HDU_PC_OUT[23] = PC_IN[23];
  assign HDU_PC_OUT[22] = PC_IN[22];
  assign HDU_PC_OUT[21] = PC_IN[21];
  assign HDU_PC_OUT[20] = PC_IN[20];
  assign HDU_PC_OUT[19] = PC_IN[19];
  assign HDU_PC_OUT[18] = PC_IN[18];
  assign HDU_PC_OUT[17] = PC_IN[17];
  assign HDU_PC_OUT[16] = PC_IN[16];
  assign HDU_PC_OUT[15] = PC_IN[15];
  assign HDU_PC_OUT[14] = PC_IN[14];
  assign HDU_PC_OUT[13] = PC_IN[13];
  assign HDU_PC_OUT[12] = PC_IN[12];
  assign HDU_PC_OUT[11] = PC_IN[11];
  assign HDU_PC_OUT[10] = PC_IN[10];
  assign HDU_PC_OUT[9] = PC_IN[9];
  assign HDU_PC_OUT[8] = PC_IN[8];
  assign HDU_PC_OUT[7] = PC_IN[7];
  assign HDU_PC_OUT[6] = PC_IN[6];
  assign HDU_PC_OUT[5] = PC_IN[5];
  assign HDU_PC_OUT[4] = PC_IN[4];
  assign HDU_PC_OUT[3] = PC_IN[3];
  assign HDU_PC_OUT[2] = PC_IN[2];
  assign HDU_PC_OUT[1] = PC_IN[1];
  assign HDU_PC_OUT[0] = PC_IN[0];

  HazardDetection_DW01_add_0 add_32 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(HDU_NPC_OUT) );
  AND3_X1 U4 ( .A1(DRAM_R), .A2(n1), .A3(RST), .ZN(Bubble) );
  OAI33_X1 U5 ( .A1(n2), .A2(n3), .A3(n4), .B1(n5), .B2(n6), .B3(n9), .ZN(n1)
         );
  XOR2_X1 U6 ( .A(ADD_WR[4]), .B(ADD_RS2[4]), .Z(n9) );
  XOR2_X1 U8 ( .A(ADD_WR[2]), .B(ADD_RS2[2]), .Z(n6) );
  NAND3_X1 U9 ( .A1(n10), .A2(n12), .A3(n13), .ZN(n5) );
  XNOR2_X1 U11 ( .A(ADD_WR[0]), .B(ADD_RS2[0]), .ZN(n13) );
  XNOR2_X1 U12 ( .A(ADD_WR[1]), .B(ADD_RS2[1]), .ZN(n12) );
  XNOR2_X1 U13 ( .A(ADD_WR[3]), .B(ADD_RS2[3]), .ZN(n10) );
  XOR2_X1 U14 ( .A(ADD_WR[4]), .B(ADD_RS1[4]), .Z(n4) );
  XOR2_X1 U15 ( .A(ADD_WR[2]), .B(ADD_RS1[2]), .Z(n3) );
  NAND3_X1 U16 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  XNOR2_X1 U17 ( .A(ADD_WR[0]), .B(ADD_RS1[0]), .ZN(n16) );
  XNOR2_X1 U18 ( .A(ADD_WR[1]), .B(ADD_RS1[1]), .ZN(n15) );
  XNOR2_X1 U19 ( .A(ADD_WR[3]), .B(ADD_RS1[3]), .ZN(n14) );
endmodule


module Datapath ( CLK, RST, INS_IN, DATA_IN, MUX_A_SEL, MUX_B_SEL, ALU_OPC, 
        ALU_OUTREG_EN, JUMP_TYPE, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE, 
        LOAD_TYPE_IN, STORE_TYPE_IN, WB_MUX_SEL, INS_OUT, IRAM_ADDR_OUT, 
        DRAM_ADDR_OUT, DATA_OUT, DRAM_R_OUT, DRAM_W_OUT, Bubble_out, 
        LOAD_TYPE_OUT, STORE_TYPE_OUT );
  input [31:0] INS_IN;
  input [31:0] DATA_IN;
  input [1:0] MUX_B_SEL;
  input [4:0] ALU_OPC;
  input [1:0] JUMP_TYPE;
  input [1:0] LOAD_TYPE_IN;
  output [31:0] INS_OUT;
  output [31:0] IRAM_ADDR_OUT;
  output [31:0] DRAM_ADDR_OUT;
  output [31:0] DATA_OUT;
  output [1:0] LOAD_TYPE_OUT;
  input CLK, RST, MUX_A_SEL, ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN,
         RF_WE, STORE_TYPE_IN, WB_MUX_SEL;
  output DRAM_R_OUT, DRAM_W_OUT, Bubble_out, STORE_TYPE_OUT;
  wire   n8, n9, n10, n11, n12, n13, n14, ZERO_FLAG_EX, RF_WE_WB, DRAM_R_MEM;
  wire   [31:0] PC_MEM_OUT;
  wire   [31:0] sig_HDU_INS_OUT;
  wire   [31:0] sig_HDU_PC_OUT;
  wire   [31:0] sig_HDU_NPC_OUT;
  wire   [31:0] PC_FETCH_OUT;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [4:0] ADD_WR_WB;
  wire   [31:0] OP_WB;
  wire   [31:0] PC_DECODE_OUT;
  wire   [31:0] A_DECODE_OUT;
  wire   [31:0] B_DECODE_OUT;
  wire   [31:0] IMM_DECODE_OUT;
  wire   [4:0] ADD_RS1_HDU;
  wire   [4:0] ADD_RS2_HDU;
  wire   [4:0] ADD_WR_DECODE_OUT;
  wire   [4:0] ADD_RS1_DECODE_OUT;
  wire   [4:0] ADD_RS2_DECODE_OUT;
  wire   [4:0] ADD_WR_MEM;
  wire   [31:0] OP_MEM;
  wire   [1:0] PC_SEL_EX;
  wire   [31:0] NPC_ABS_EX;
  wire   [31:0] NPC_REL_EX;
  wire   [31:0] ALU_RES_EX;
  wire   [31:0] B_EX_OUT;
  wire   [4:0] ADD_WR_EX_OUT;
  wire   [31:0] DATA_MEM_OUT;
  wire   [31:0] ALU_RES_MEM;
  wire   [4:0] ADD_WR_MEM_OUT;

  Fetch FetchStage ( .CLK(CLK), .RST(RST), .ZERO_FLAG(ZERO_FLAG_EX), .PC_EXT(
        PC_MEM_OUT), .INS_IN(INS_IN), .Bubble_in(Bubble_out), .HDU_INS_IN(
        sig_HDU_INS_OUT), .HDU_PC_IN(sig_HDU_PC_OUT), .HDU_NPC_IN(
        sig_HDU_NPC_OUT), .PC_OUT(PC_FETCH_OUT), .ADDR_OUT(IRAM_ADDR_OUT), 
        .NPC_OUT(NPC_FETCH_OUT), .INS_OUT({n8, n9, n10, n11, n12, n13, 
        INS_OUT[25:0]}) );
  Decode DecodeStage ( .CLK(CLK), .RST(RST), .Bubble(Bubble_out), .RF_WE(
        RF_WE_WB), .ZERO_FLAG(ZERO_FLAG_EX), .PC_IN(PC_FETCH_OUT), .INS_IN({n8, 
        n9, n10, n11, n12, n13, INS_OUT[25:0]}), .ADD_WR(ADD_WR_WB), 
        .DATA_WR_IN(OP_WB), .PC_OUT(PC_DECODE_OUT), .A_OUT(A_DECODE_OUT), 
        .B_OUT(B_DECODE_OUT), .IMM_OUT(IMM_DECODE_OUT), .ADD_RS1_HDU(
        ADD_RS1_HDU), .ADD_RS2_HDU(ADD_RS2_HDU), .ADD_WR_OUT(ADD_WR_DECODE_OUT), .ADD_RS1_OUT(ADD_RS1_DECODE_OUT), .ADD_RS2_OUT(ADD_RS2_DECODE_OUT) );
  Execute ExecuteStage ( .CLK(CLK), .RST(RST), .MUX_A_SEL(MUX_A_SEL), 
        .MUX_B_SEL(MUX_B_SEL), .ALU_OPC(ALU_OPC), .ALU_OUTREG_EN(ALU_OUTREG_EN), .JUMP_TYPE(JUMP_TYPE), .PC_IN(PC_DECODE_OUT), .A_IN(A_DECODE_OUT), .B_IN(
        B_DECODE_OUT), .IMM_IN(IMM_DECODE_OUT), .ADD_WR_IN(ADD_WR_DECODE_OUT), 
        .ADD_RS1_IN(ADD_RS1_DECODE_OUT), .ADD_RS2_IN(ADD_RS2_DECODE_OUT), 
        .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_WB(ADD_WR_WB), .RF_WE_MEM(RF_WE), 
        .RF_WE_WB(RF_WE_WB), .OP_MEM(OP_MEM), .OP_WB(OP_WB), .PC_SEL(PC_SEL_EX), .ZERO_FLAG(ZERO_FLAG_EX), .NPC_ABS(NPC_ABS_EX), .NPC_REL(NPC_REL_EX), 
        .ALU_RES(ALU_RES_EX), .B_OUT(B_EX_OUT), .ADD_WR_OUT(ADD_WR_EX_OUT) );
  ff_0 DRAM_R_ff ( .D(DRAM_R_IN), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DRAM_R_MEM) );
  Memory MemoryStage ( .CLK(CLK), .RST(RST), .MEM_EN_IN(MEM_EN_IN), 
        .DRAM_R_IN(DRAM_R_MEM), .DRAM_W_IN(DRAM_W_IN), .PC_SEL(PC_SEL_EX), 
        .NPC_IN(NPC_FETCH_OUT), .NPC_ABS(NPC_ABS_EX), .NPC_REL(NPC_REL_EX), 
        .ALU_RES_IN(ALU_RES_EX), .B_IN(B_EX_OUT), .ADD_WR_IN(ADD_WR_EX_OUT), 
        .DRAM_DATA_IN(DATA_IN), .LOAD_TYPE_IN(LOAD_TYPE_IN), .STORE_TYPE_IN(
        STORE_TYPE_IN), .PC_OUT(PC_MEM_OUT), .DRAM_R_OUT(DRAM_R_OUT), 
        .DRAM_W_OUT(DRAM_W_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DRAM_DATA_OUT(DATA_OUT), .DATA_OUT(DATA_MEM_OUT), .ALU_RES_OUT(
        ALU_RES_MEM), .OP_MEM(OP_MEM), .ADD_WR_MEM(ADD_WR_MEM), .ADD_WR_OUT(
        ADD_WR_MEM_OUT), .LOAD_TYPE_OUT(LOAD_TYPE_OUT), .STORE_TYPE_OUT(
        STORE_TYPE_OUT) );
  ff_2 RF_WE_ff ( .D(RF_WE), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(RF_WE_WB) );
  Writeback WritebackStage ( .WB_MUX_SEL(WB_MUX_SEL), .DATA_IN(DATA_MEM_OUT), 
        .ALU_RES_IN(ALU_RES_MEM), .ADD_WR_IN(ADD_WR_MEM_OUT), .DATA_OUT(OP_WB), 
        .ADD_WR_OUT(ADD_WR_WB) );
  HazardDetection HDU ( .RST(RST), .ADD_RS1(ADD_RS1_HDU), .ADD_RS2(ADD_RS2_HDU), .ADD_WR(ADD_WR_DECODE_OUT), .DRAM_R(DRAM_R_IN), .INS_IN(INS_OUT), .PC_IN(
        PC_FETCH_OUT), .Bubble(n14), .HDU_INS_OUT(sig_HDU_INS_OUT), 
        .HDU_PC_OUT(sig_HDU_PC_OUT), .HDU_NPC_OUT(sig_HDU_NPC_OUT) );
  BUF_X1 U2 ( .A(n14), .Z(Bubble_out) );
  CLKBUF_X1 U3 ( .A(n10), .Z(INS_OUT[29]) );
  CLKBUF_X1 U4 ( .A(n12), .Z(INS_OUT[27]) );
  CLKBUF_X1 U5 ( .A(n13), .Z(INS_OUT[26]) );
  CLKBUF_X1 U6 ( .A(n9), .Z(INS_OUT[30]) );
  CLKBUF_X1 U7 ( .A(n11), .Z(INS_OUT[28]) );
  CLKBUF_X1 U8 ( .A(n8), .Z(INS_OUT[31]) );
endmodule


module hardwired_cu_NBIT32 ( MUX_A_SEL, MUX_B_SEL, ALU_OPC, ALU_OUTREG_EN, 
        DRAM_R_IN, JUMP_TYPE, MEM_EN_IN, DRAM_W_IN, RF_WE, LOAD_TYPE_IN, 
        STORE_TYPE_IN, WB_MUX_SEL, INS_IN, Bubble, Clk, Rst );
  output [1:0] MUX_B_SEL;
  output [4:0] ALU_OPC;
  output [1:0] JUMP_TYPE;
  output [1:0] LOAD_TYPE_IN;
  input [31:0] INS_IN;
  input Bubble, Clk, Rst;
  output MUX_A_SEL, ALU_OUTREG_EN, DRAM_R_IN, MEM_EN_IN, DRAM_W_IN, RF_WE,
         STORE_TYPE_IN, WB_MUX_SEL;
  wire   n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28;
  wire   [4:0] AluOP_E;
  assign MUX_A_SEL = 1'b0;
  assign MUX_B_SEL[1] = 1'b0;
  assign MUX_B_SEL[0] = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign DRAM_R_IN = 1'b0;
  assign JUMP_TYPE[1] = 1'b0;
  assign JUMP_TYPE[0] = 1'b0;
  assign MEM_EN_IN = 1'b0;
  assign DRAM_W_IN = 1'b0;
  assign RF_WE = 1'b0;
  assign LOAD_TYPE_IN[1] = 1'b0;
  assign LOAD_TYPE_IN[0] = 1'b0;
  assign STORE_TYPE_IN = 1'b0;
  assign WB_MUX_SEL = 1'b0;

  DFFR_X1 ALU_OPC_reg_0_ ( .D(AluOP_E[0]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[0])
         );
  NAND3_X1 U126 ( .A1(INS_IN[1]), .A2(n25), .A3(INS_IN[0]), .ZN(n65) );
  NAND3_X1 U127 ( .A1(n87), .A2(n64), .A3(n88), .ZN(n51) );
  XOR2_X1 U128 ( .A(n28), .B(INS_IN[1]), .Z(n91) );
  NAND3_X1 U129 ( .A1(n92), .A2(n27), .A3(INS_IN[0]), .ZN(n37) );
  NAND3_X1 U130 ( .A1(n10), .A2(n7), .A3(n33), .ZN(n103) );
  NAND3_X1 U131 ( .A1(n28), .A2(n27), .A3(n92), .ZN(n39) );
  NAND3_X1 U132 ( .A1(n110), .A2(n25), .A3(INS_IN[1]), .ZN(n38) );
  NAND3_X1 U133 ( .A1(n26), .A2(n27), .A3(n53), .ZN(n106) );
  NAND3_X1 U134 ( .A1(INS_IN[1]), .A2(n28), .A3(n92), .ZN(n43) );
  NAND3_X1 U135 ( .A1(n23), .A2(n21), .A3(n113), .ZN(n112) );
  DFFR_X1 ALU_OPC_reg_3_ ( .D(AluOP_E[3]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[3])
         );
  DFFR_X1 ALU_OPC_reg_1_ ( .D(AluOP_E[1]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[1])
         );
  DFFR_X1 ALU_OPC_reg_4_ ( .D(AluOP_E[4]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[4])
         );
  DFFR_X1 ALU_OPC_reg_2_ ( .D(AluOP_E[2]), .CK(Clk), .RN(Rst), .Q(ALU_OPC[2])
         );
  INV_X1 U17 ( .A(n79), .ZN(n4) );
  NAND2_X1 U18 ( .A1(n82), .A2(n66), .ZN(n73) );
  INV_X1 U19 ( .A(n82), .ZN(n5) );
  INV_X1 U20 ( .A(n66), .ZN(n2) );
  INV_X1 U21 ( .A(n34), .ZN(n13) );
  NOR3_X1 U22 ( .A1(n33), .A2(n99), .A3(n11), .ZN(n81) );
  INV_X1 U23 ( .A(n77), .ZN(n11) );
  NAND2_X1 U24 ( .A1(n70), .A2(n8), .ZN(n79) );
  NAND2_X1 U25 ( .A1(n70), .A2(n9), .ZN(n82) );
  NAND2_X1 U26 ( .A1(n68), .A2(n69), .ZN(n54) );
  OAI21_X1 U27 ( .B1(n100), .B2(n75), .A(n101), .ZN(n95) );
  NOR3_X1 U28 ( .A1(n102), .A2(n4), .A3(n46), .ZN(n100) );
  OAI21_X1 U29 ( .B1(n14), .B2(n57), .A(n73), .ZN(n101) );
  OAI21_X1 U30 ( .B1(n3), .B2(n60), .A(n103), .ZN(n102) );
  AND4_X1 U31 ( .A1(n70), .A2(n57), .A3(n10), .A4(n7), .ZN(n35) );
  NAND2_X1 U32 ( .A1(n75), .A2(n59), .ZN(n34) );
  NAND2_X1 U33 ( .A1(n9), .A2(n74), .ZN(n66) );
  INV_X1 U34 ( .A(n60), .ZN(n9) );
  INV_X1 U35 ( .A(n75), .ZN(n12) );
  INV_X1 U36 ( .A(n59), .ZN(n14) );
  OAI221_X1 U37 ( .B1(n78), .B2(n79), .C1(n66), .C2(n11), .A(n80), .ZN(n67) );
  NOR3_X1 U38 ( .A1(n77), .A2(n57), .A3(n12), .ZN(n78) );
  NOR2_X1 U39 ( .A1(n48), .A2(n81), .ZN(n80) );
  AND3_X1 U40 ( .A1(n8), .A2(n74), .A3(n57), .ZN(n32) );
  AND3_X1 U41 ( .A1(n8), .A2(n74), .A3(n77), .ZN(n48) );
  INV_X1 U42 ( .A(n105), .ZN(n1) );
  AOI21_X1 U43 ( .B1(n57), .B2(n46), .A(n81), .ZN(n105) );
  INV_X1 U44 ( .A(n99), .ZN(n8) );
  INV_X1 U45 ( .A(n51), .ZN(n17) );
  AOI21_X1 U46 ( .B1(n44), .B2(n45), .A(Bubble), .ZN(AluOP_E[3]) );
  AOI211_X1 U47 ( .C1(n14), .C2(n4), .A(n54), .B(n1), .ZN(n44) );
  AOI221_X1 U48 ( .B1(n46), .B2(n34), .C1(n35), .C2(n47), .A(n48), .ZN(n45) );
  OAI21_X1 U49 ( .B1(n49), .B2(n50), .A(n17), .ZN(n47) );
  AOI21_X1 U50 ( .B1(n93), .B2(n94), .A(Bubble), .ZN(AluOP_E[0]) );
  NOR3_X1 U51 ( .A1(n95), .A2(n6), .A3(n96), .ZN(n94) );
  AOI221_X1 U52 ( .B1(n35), .B2(n104), .C1(n77), .C2(n4), .A(n1), .ZN(n93) );
  INV_X1 U53 ( .A(n68), .ZN(n6) );
  AOI22_X1 U54 ( .A1(n98), .A2(n77), .B1(n57), .B2(n99), .ZN(n97) );
  NAND2_X1 U55 ( .A1(n52), .A2(n89), .ZN(n83) );
  AOI21_X1 U56 ( .B1(n29), .B2(n30), .A(Bubble), .ZN(AluOP_E[4]) );
  AOI211_X1 U57 ( .C1(n31), .C2(n9), .A(n2), .B(n32), .ZN(n30) );
  AOI22_X1 U58 ( .A1(n35), .A2(n36), .B1(n12), .B2(n4), .ZN(n29) );
  NOR2_X1 U59 ( .A1(n13), .A2(n33), .ZN(n31) );
  OAI21_X1 U60 ( .B1(n52), .B2(n41), .A(n27), .ZN(n90) );
  NAND4_X1 U61 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n36) );
  AOI21_X1 U62 ( .B1(n41), .B2(n42), .A(n20), .ZN(n40) );
  INV_X1 U63 ( .A(n43), .ZN(n20) );
  AOI21_X1 U64 ( .B1(n55), .B2(n56), .A(Bubble), .ZN(AluOP_E[2]) );
  AOI211_X1 U65 ( .C1(n5), .C2(n12), .A(n67), .B(n54), .ZN(n55) );
  AOI221_X1 U66 ( .B1(n2), .B2(n57), .C1(n35), .C2(n16), .A(n58), .ZN(n56) );
  NOR3_X1 U67 ( .A1(n59), .A2(n33), .A3(n60), .ZN(n58) );
  NAND2_X1 U68 ( .A1(n89), .A2(n110), .ZN(n87) );
  NAND2_X1 U69 ( .A1(n89), .A2(n41), .ZN(n64) );
  AOI21_X1 U70 ( .B1(n71), .B2(n72), .A(Bubble), .ZN(AluOP_E[1]) );
  AOI221_X1 U71 ( .B1(n46), .B2(n34), .C1(n14), .C2(n73), .A(n32), .ZN(n72) );
  AOI221_X1 U72 ( .B1(n35), .B2(n76), .C1(n5), .C2(n77), .A(n67), .ZN(n71) );
  NAND4_X1 U73 ( .A1(n43), .A2(n37), .A3(n83), .A4(n84), .ZN(n76) );
  INV_X1 U74 ( .A(n53), .ZN(n19) );
  INV_X1 U75 ( .A(n38), .ZN(n18) );
  AND2_X1 U76 ( .A1(n41), .A2(n25), .ZN(n92) );
  INV_X1 U77 ( .A(n50), .ZN(n26) );
  NOR3_X1 U78 ( .A1(n22), .A2(INS_IN[3]), .A3(n112), .ZN(n52) );
  NOR3_X1 U79 ( .A1(n22), .A2(n24), .A3(n112), .ZN(n41) );
  INV_X1 U80 ( .A(INS_IN[3]), .ZN(n24) );
  NOR3_X1 U81 ( .A1(INS_IN[3]), .A2(INS_IN[5]), .A3(n112), .ZN(n53) );
  NOR3_X1 U82 ( .A1(n28), .A2(INS_IN[1]), .A3(n25), .ZN(n89) );
  NOR4_X1 U83 ( .A1(INS_IN[7]), .A2(INS_IN[10]), .A3(INS_IN[9]), .A4(INS_IN[8]), .ZN(n113) );
  AOI221_X1 U84 ( .B1(n85), .B2(n52), .C1(n26), .C2(n86), .A(n51), .ZN(n84) );
  NOR2_X1 U85 ( .A1(INS_IN[2]), .A2(n91), .ZN(n85) );
  OAI21_X1 U86 ( .B1(n27), .B2(n19), .A(n90), .ZN(n86) );
  NAND4_X1 U87 ( .A1(n88), .A2(n43), .A3(n106), .A4(n107), .ZN(n104) );
  AOI221_X1 U88 ( .B1(n108), .B2(n52), .C1(n18), .C2(INS_IN[0]), .A(n62), .ZN(
        n107) );
  NOR2_X1 U89 ( .A1(INS_IN[2]), .A2(INS_IN[0]), .ZN(n108) );
  OAI21_X1 U90 ( .B1(INS_IN[1]), .B2(n50), .A(n65), .ZN(n42) );
  NAND4_X1 U91 ( .A1(n53), .A2(INS_IN[2]), .A3(INS_IN[0]), .A4(INS_IN[1]), 
        .ZN(n88) );
  NAND2_X1 U92 ( .A1(INS_IN[2]), .A2(n28), .ZN(n50) );
  INV_X1 U93 ( .A(INS_IN[1]), .ZN(n27) );
  AOI21_X1 U94 ( .B1(n52), .B2(INS_IN[1]), .A(n53), .ZN(n49) );
  NAND4_X1 U95 ( .A1(n109), .A2(n83), .A3(n87), .A4(n39), .ZN(n62) );
  NAND4_X1 U96 ( .A1(INS_IN[3]), .A2(n22), .A3(INS_IN[1]), .A4(n111), .ZN(n109) );
  NOR2_X1 U97 ( .A1(n112), .A2(n50), .ZN(n111) );
  INV_X1 U98 ( .A(INS_IN[0]), .ZN(n28) );
  INV_X1 U99 ( .A(INS_IN[5]), .ZN(n22) );
  INV_X1 U100 ( .A(INS_IN[2]), .ZN(n25) );
  AND4_X1 U101 ( .A1(n113), .A2(n21), .A3(INS_IN[3]), .A4(n114), .ZN(n110) );
  NOR2_X1 U102 ( .A1(n23), .A2(n22), .ZN(n114) );
  INV_X1 U103 ( .A(INS_IN[4]), .ZN(n23) );
  INV_X1 U104 ( .A(INS_IN[6]), .ZN(n21) );
  INV_X1 U105 ( .A(n61), .ZN(n16) );
  AOI211_X1 U106 ( .C1(n42), .C2(n52), .A(n62), .B(n63), .ZN(n61) );
  OAI211_X1 U107 ( .C1(n38), .C2(INS_IN[0]), .A(n37), .B(n64), .ZN(n63) );
  NOR2_X1 U108 ( .A1(INS_IN[29]), .A2(n10), .ZN(n98) );
  INV_X1 U109 ( .A(INS_IN[29]), .ZN(n7) );
  NAND2_X1 U110 ( .A1(INS_IN[29]), .A2(n10), .ZN(n60) );
  INV_X1 U111 ( .A(INS_IN[26]), .ZN(n15) );
  NOR3_X1 U112 ( .A1(n3), .A2(INS_IN[30]), .A3(n97), .ZN(n96) );
  AND2_X1 U113 ( .A1(INS_IN[30]), .A2(n3), .ZN(n74) );
  NAND2_X1 U114 ( .A1(INS_IN[27]), .A2(n15), .ZN(n59) );
  NAND2_X1 U115 ( .A1(INS_IN[26]), .A2(INS_IN[27]), .ZN(n75) );
  NOR2_X1 U116 ( .A1(n15), .A2(INS_IN[27]), .ZN(n77) );
  NOR2_X1 U117 ( .A1(INS_IN[27]), .A2(INS_IN[26]), .ZN(n57) );
  NAND4_X1 U118 ( .A1(n70), .A2(n57), .A3(INS_IN[28]), .A4(n7), .ZN(n69) );
  NAND4_X1 U119 ( .A1(n77), .A2(n70), .A3(INS_IN[28]), .A4(n7), .ZN(n68) );
  AND3_X1 U120 ( .A1(INS_IN[28]), .A2(n7), .A3(n74), .ZN(n46) );
  NAND2_X1 U121 ( .A1(INS_IN[29]), .A2(INS_IN[28]), .ZN(n99) );
  INV_X1 U122 ( .A(INS_IN[28]), .ZN(n10) );
  NAND2_X1 U123 ( .A1(INS_IN[31]), .A2(INS_IN[30]), .ZN(n33) );
  NOR2_X1 U124 ( .A1(INS_IN[31]), .A2(INS_IN[30]), .ZN(n70) );
  INV_X1 U125 ( .A(INS_IN[31]), .ZN(n3) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   DRAM_R_OUT, DRAM_W_OUT, Bubble, STORE_TYPE_OUT,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6;
  wire   [31:0] INS_IN;
  wire   [31:0] DATA_IN;
  wire   [1:0] MUX_B_SEL;
  wire   [4:0] ALU_OPC;
  wire   [1:0] JUMP_TYPE;
  wire   [1:0] LOAD_TYPE_IN;
  wire   [31:0] INST;
  wire   [31:0] IRAM_ADDR_OUT;
  wire   [31:0] DRAM_ADDR_OUT;
  wire   [31:0] DATA_OUT;
  wire   [1:0] LOAD_TYPE_OUT;

  Datapath DP ( .CLK(Clk), .RST(Rst), .INS_IN(INS_IN), .DATA_IN(DATA_IN), 
        .MUX_A_SEL(1'b0), .MUX_B_SEL({1'b0, 1'b0}), .ALU_OPC(ALU_OPC), 
        .ALU_OUTREG_EN(1'b0), .JUMP_TYPE({1'b0, 1'b0}), .DRAM_R_IN(1'b0), 
        .MEM_EN_IN(1'b0), .DRAM_W_IN(1'b0), .RF_WE(1'b0), .LOAD_TYPE_IN({1'b0, 
        1'b0}), .STORE_TYPE_IN(1'b0), .WB_MUX_SEL(1'b0), .INS_OUT(INST), 
        .IRAM_ADDR_OUT(IRAM_ADDR_OUT), .DRAM_ADDR_OUT(DRAM_ADDR_OUT), 
        .DATA_OUT(DATA_OUT), .DRAM_R_OUT(DRAM_R_OUT), .DRAM_W_OUT(DRAM_W_OUT), 
        .Bubble_out(Bubble), .LOAD_TYPE_OUT(LOAD_TYPE_OUT), .STORE_TYPE_OUT(
        STORE_TYPE_OUT) );
  hardwired_cu_NBIT32 CU ( .MUX_B_SEL({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .ALU_OPC(ALU_OPC), .JUMP_TYPE({
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}), .LOAD_TYPE_IN({
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}), .INS_IN(INST), 
        .Bubble(Bubble), .Clk(Clk), .Rst(Rst) );
  IRAM IRAM_I ( .Rst(Rst), .Addr(IRAM_ADDR_OUT), .Iout(INS_IN) );
  DRAM DRAM_I ( .Clk(Clk), .Rst(Rst), .ADDR_IN(DRAM_ADDR_OUT), .DATA_IN(
        DATA_OUT), .LOAD_TYPE(LOAD_TYPE_OUT), .STORE_TYPE(STORE_TYPE_OUT), 
        .DRAM_W(DRAM_W_OUT), .DRAM_R(DRAM_R_OUT), .DATA_OUT(DATA_IN) );
endmodule

