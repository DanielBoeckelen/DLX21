library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use work.constants.all;

entity tb_comparator is
end entity;

architecture test of tb_comparator is

component comparator is
	generic(NBIT : integer);
	port(     A     : in std_logic_vector(NBIT-1 downto 0);
		  B     : in std_logic_vector(NBIT-1 downto 0);
		  OPSel : in integer range 0 to 5;
		  RES   : out std_logic_vector(NBIT-1 downto 0));
end component;

  constant tb_period : time := 10ns;

   signal A : std_logic_vector(NBIT-1 downto 0);
   signal B : std_logic_vector(NBIT-1 downto 0);
   signal OPSel : integer range 0 to 5;
   signal RES   : std_logic_vector(NBIT-1 downto 0);

begin

  DUT : comparator
    generic map (NBIT => 32)
    port map(
                 A => A,
                 B => B,
                 OPSel => OPSel,
                 RES => RES
                );

  stimuli : process

                procedure apply_stimuli (
                        constant A_val : in integer;
                        constant B_val : in integer;
                        constant OPSel_val : in integer range 0 to 5;
                        
                        signal A : out std_logic_vector(NBIT-1 downto 0);
                        signal B : out std_logic_vector(NBIT-1 downto 0);
                        signal OPSel : out integer range 0 to 5) is
                begin
                       A <= conv_std_logic_vector(A_val, NBIT); --integer
                       B <= conv_std_logic_vector(B_val, NBIT); --integer
                       OPSel <= OPSel_val;
	
                        --A <= A_val; --hex
                        --B <= B_val; --hex
                       
                        wait for tb_period;
                       
                end apply_stimuli;
  begin

   --apply_stimuli(input values, signals);

 -- a < b
  for i in 0 to 5 loop
    
    apply_stimuli(0, 1, i, A, B, OPSel);
    
  end loop;

 -- a = b
 for i in 0 to 5 loop
    
    apply_stimuli(7, 7, i, A, B, OPSel);
    
 end loop;

-- a > b  
for i in 0 to 5 loop
    
   apply_stimuli(26, 21, i, A, B, OPSel);
    
end loop;
  
  end process;

end test;
