library verilog;
use verilog.vl_types.all;
entity DLX is
    port(
        Clk             : in     vl_logic;
        Rst             : in     vl_logic
    );
end DLX;
