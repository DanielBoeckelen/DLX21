library verilog;
use verilog.vl_types.all;
entity Gblock_1 is
    port(
        Pik             : in     vl_logic;
        Gik             : in     vl_logic;
        Gk_1j           : in     vl_logic;
        Gij             : out    vl_logic
    );
end Gblock_1;
