ms21.21@localhost.localdomain.8325:1614348791